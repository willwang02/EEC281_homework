`timescale 10ps/1ps

module prob1_2 (
    clk,
    theta,
    out
);
    input clk;
    input [11:0] theta;
    output reg [15:0] out;
    reg [16:0] out_r;
    reg [16:0] lvalue_r, rvalue_r;
    reg even;
    always @(posedge clk) begin
        case(theta >> 1)
            11'b00000000000: begin lvalue_r <= 16'b0000000000000000; rvalue_r <= 16'b0000000000001101;end
            11'b00000000001: begin lvalue_r <= 16'b0000000000001101; rvalue_r <= 16'b0000000000011001;end
            11'b00000000010: begin lvalue_r <= 16'b0000000000011001; rvalue_r <= 16'b0000000000100110;end
            11'b00000000011: begin lvalue_r <= 16'b0000000000100110; rvalue_r <= 16'b0000000000110010;end
            11'b00000000100: begin lvalue_r <= 16'b0000000000110010; rvalue_r <= 16'b0000000000111111;end
            11'b00000000101: begin lvalue_r <= 16'b0000000000111111; rvalue_r <= 16'b0000000001001011;end
            11'b00000000110: begin lvalue_r <= 16'b0000000001001011; rvalue_r <= 16'b0000000001011000;end
            11'b00000000111: begin lvalue_r <= 16'b0000000001011000; rvalue_r <= 16'b0000000001100101;end
            11'b00000001000: begin lvalue_r <= 16'b0000000001100101; rvalue_r <= 16'b0000000001110001;end
            11'b00000001001: begin lvalue_r <= 16'b0000000001110001; rvalue_r <= 16'b0000000001111110;end
            11'b00000001010: begin lvalue_r <= 16'b0000000001111110; rvalue_r <= 16'b0000000010001010;end
            11'b00000001011: begin lvalue_r <= 16'b0000000010001010; rvalue_r <= 16'b0000000010010111;end
            11'b00000001100: begin lvalue_r <= 16'b0000000010010111; rvalue_r <= 16'b0000000010100011;end
            11'b00000001101: begin lvalue_r <= 16'b0000000010100011; rvalue_r <= 16'b0000000010110000;end
            11'b00000001110: begin lvalue_r <= 16'b0000000010110000; rvalue_r <= 16'b0000000010111100;end
            11'b00000001111: begin lvalue_r <= 16'b0000000010111100; rvalue_r <= 16'b0000000011001001;end
            11'b00000010000: begin lvalue_r <= 16'b0000000011001001; rvalue_r <= 16'b0000000011010110;end
            11'b00000010001: begin lvalue_r <= 16'b0000000011010110; rvalue_r <= 16'b0000000011100010;end
            11'b00000010010: begin lvalue_r <= 16'b0000000011100010; rvalue_r <= 16'b0000000011101111;end
            11'b00000010011: begin lvalue_r <= 16'b0000000011101111; rvalue_r <= 16'b0000000011111011;end
            11'b00000010100: begin lvalue_r <= 16'b0000000011111011; rvalue_r <= 16'b0000000100001000;end
            11'b00000010101: begin lvalue_r <= 16'b0000000100001000; rvalue_r <= 16'b0000000100010100;end
            11'b00000010110: begin lvalue_r <= 16'b0000000100010100; rvalue_r <= 16'b0000000100100001;end
            11'b00000010111: begin lvalue_r <= 16'b0000000100100001; rvalue_r <= 16'b0000000100101110;end
            11'b00000011000: begin lvalue_r <= 16'b0000000100101110; rvalue_r <= 16'b0000000100111010;end
            11'b00000011001: begin lvalue_r <= 16'b0000000100111010; rvalue_r <= 16'b0000000101000111;end
            11'b00000011010: begin lvalue_r <= 16'b0000000101000111; rvalue_r <= 16'b0000000101010011;end
            11'b00000011011: begin lvalue_r <= 16'b0000000101010011; rvalue_r <= 16'b0000000101100000;end
            11'b00000011100: begin lvalue_r <= 16'b0000000101100000; rvalue_r <= 16'b0000000101101100;end
            11'b00000011101: begin lvalue_r <= 16'b0000000101101100; rvalue_r <= 16'b0000000101111001;end
            11'b00000011110: begin lvalue_r <= 16'b0000000101111001; rvalue_r <= 16'b0000000110000110;end
            11'b00000011111: begin lvalue_r <= 16'b0000000110000110; rvalue_r <= 16'b0000000110010010;end
            11'b00000100000: begin lvalue_r <= 16'b0000000110010010; rvalue_r <= 16'b0000000110011111;end
            11'b00000100001: begin lvalue_r <= 16'b0000000110011111; rvalue_r <= 16'b0000000110101011;end
            11'b00000100010: begin lvalue_r <= 16'b0000000110101011; rvalue_r <= 16'b0000000110111000;end
            11'b00000100011: begin lvalue_r <= 16'b0000000110111000; rvalue_r <= 16'b0000000111000100;end
            11'b00000100100: begin lvalue_r <= 16'b0000000111000100; rvalue_r <= 16'b0000000111010001;end
            11'b00000100101: begin lvalue_r <= 16'b0000000111010001; rvalue_r <= 16'b0000000111011110;end
            11'b00000100110: begin lvalue_r <= 16'b0000000111011110; rvalue_r <= 16'b0000000111101010;end
            11'b00000100111: begin lvalue_r <= 16'b0000000111101010; rvalue_r <= 16'b0000000111110111;end
            11'b00000101000: begin lvalue_r <= 16'b0000000111110111; rvalue_r <= 16'b0000001000000011;end
            11'b00000101001: begin lvalue_r <= 16'b0000001000000011; rvalue_r <= 16'b0000001000010000;end
            11'b00000101010: begin lvalue_r <= 16'b0000001000010000; rvalue_r <= 16'b0000001000011100;end
            11'b00000101011: begin lvalue_r <= 16'b0000001000011100; rvalue_r <= 16'b0000001000101001;end
            11'b00000101100: begin lvalue_r <= 16'b0000001000101001; rvalue_r <= 16'b0000001000110110;end
            11'b00000101101: begin lvalue_r <= 16'b0000001000110110; rvalue_r <= 16'b0000001001000010;end
            11'b00000101110: begin lvalue_r <= 16'b0000001001000010; rvalue_r <= 16'b0000001001001111;end
            11'b00000101111: begin lvalue_r <= 16'b0000001001001111; rvalue_r <= 16'b0000001001011011;end
            11'b00000110000: begin lvalue_r <= 16'b0000001001011011; rvalue_r <= 16'b0000001001101000;end
            11'b00000110001: begin lvalue_r <= 16'b0000001001101000; rvalue_r <= 16'b0000001001110100;end
            11'b00000110010: begin lvalue_r <= 16'b0000001001110100; rvalue_r <= 16'b0000001010000001;end
            11'b00000110011: begin lvalue_r <= 16'b0000001010000001; rvalue_r <= 16'b0000001010001110;end
            11'b00000110100: begin lvalue_r <= 16'b0000001010001110; rvalue_r <= 16'b0000001010011010;end
            11'b00000110101: begin lvalue_r <= 16'b0000001010011010; rvalue_r <= 16'b0000001010100111;end
            11'b00000110110: begin lvalue_r <= 16'b0000001010100111; rvalue_r <= 16'b0000001010110011;end
            11'b00000110111: begin lvalue_r <= 16'b0000001010110011; rvalue_r <= 16'b0000001011000000;end
            11'b00000111000: begin lvalue_r <= 16'b0000001011000000; rvalue_r <= 16'b0000001011001100;end
            11'b00000111001: begin lvalue_r <= 16'b0000001011001100; rvalue_r <= 16'b0000001011011001;end
            11'b00000111010: begin lvalue_r <= 16'b0000001011011001; rvalue_r <= 16'b0000001011100110;end
            11'b00000111011: begin lvalue_r <= 16'b0000001011100110; rvalue_r <= 16'b0000001011110010;end
            11'b00000111100: begin lvalue_r <= 16'b0000001011110010; rvalue_r <= 16'b0000001011111111;end
            11'b00000111101: begin lvalue_r <= 16'b0000001011111111; rvalue_r <= 16'b0000001100001011;end
            11'b00000111110: begin lvalue_r <= 16'b0000001100001011; rvalue_r <= 16'b0000001100011000;end
            11'b00000111111: begin lvalue_r <= 16'b0000001100011000; rvalue_r <= 16'b0000001100100100;end
            11'b00001000000: begin lvalue_r <= 16'b0000001100100100; rvalue_r <= 16'b0000001100110001;end
            11'b00001000001: begin lvalue_r <= 16'b0000001100110001; rvalue_r <= 16'b0000001100111110;end
            11'b00001000010: begin lvalue_r <= 16'b0000001100111110; rvalue_r <= 16'b0000001101001010;end
            11'b00001000011: begin lvalue_r <= 16'b0000001101001010; rvalue_r <= 16'b0000001101010111;end
            11'b00001000100: begin lvalue_r <= 16'b0000001101010111; rvalue_r <= 16'b0000001101100011;end
            11'b00001000101: begin lvalue_r <= 16'b0000001101100011; rvalue_r <= 16'b0000001101110000;end
            11'b00001000110: begin lvalue_r <= 16'b0000001101110000; rvalue_r <= 16'b0000001101111100;end
            11'b00001000111: begin lvalue_r <= 16'b0000001101111100; rvalue_r <= 16'b0000001110001001;end
            11'b00001001000: begin lvalue_r <= 16'b0000001110001001; rvalue_r <= 16'b0000001110010110;end
            11'b00001001001: begin lvalue_r <= 16'b0000001110010110; rvalue_r <= 16'b0000001110100010;end
            11'b00001001010: begin lvalue_r <= 16'b0000001110100010; rvalue_r <= 16'b0000001110101111;end
            11'b00001001011: begin lvalue_r <= 16'b0000001110101111; rvalue_r <= 16'b0000001110111011;end
            11'b00001001100: begin lvalue_r <= 16'b0000001110111011; rvalue_r <= 16'b0000001111001000;end
            11'b00001001101: begin lvalue_r <= 16'b0000001111001000; rvalue_r <= 16'b0000001111010100;end
            11'b00001001110: begin lvalue_r <= 16'b0000001111010100; rvalue_r <= 16'b0000001111100001;end
            11'b00001001111: begin lvalue_r <= 16'b0000001111100001; rvalue_r <= 16'b0000001111101110;end
            11'b00001010000: begin lvalue_r <= 16'b0000001111101110; rvalue_r <= 16'b0000001111111010;end
            11'b00001010001: begin lvalue_r <= 16'b0000001111111010; rvalue_r <= 16'b0000010000000111;end
            11'b00001010010: begin lvalue_r <= 16'b0000010000000111; rvalue_r <= 16'b0000010000010011;end
            11'b00001010011: begin lvalue_r <= 16'b0000010000010011; rvalue_r <= 16'b0000010000100000;end
            11'b00001010100: begin lvalue_r <= 16'b0000010000100000; rvalue_r <= 16'b0000010000101101;end
            11'b00001010101: begin lvalue_r <= 16'b0000010000101101; rvalue_r <= 16'b0000010000111001;end
            11'b00001010110: begin lvalue_r <= 16'b0000010000111001; rvalue_r <= 16'b0000010001000110;end
            11'b00001010111: begin lvalue_r <= 16'b0000010001000110; rvalue_r <= 16'b0000010001010010;end
            11'b00001011000: begin lvalue_r <= 16'b0000010001010010; rvalue_r <= 16'b0000010001011111;end
            11'b00001011001: begin lvalue_r <= 16'b0000010001011111; rvalue_r <= 16'b0000010001101011;end
            11'b00001011010: begin lvalue_r <= 16'b0000010001101011; rvalue_r <= 16'b0000010001111000;end
            11'b00001011011: begin lvalue_r <= 16'b0000010001111000; rvalue_r <= 16'b0000010010000101;end
            11'b00001011100: begin lvalue_r <= 16'b0000010010000101; rvalue_r <= 16'b0000010010010001;end
            11'b00001011101: begin lvalue_r <= 16'b0000010010010001; rvalue_r <= 16'b0000010010011110;end
            11'b00001011110: begin lvalue_r <= 16'b0000010010011110; rvalue_r <= 16'b0000010010101010;end
            11'b00001011111: begin lvalue_r <= 16'b0000010010101010; rvalue_r <= 16'b0000010010110111;end
            11'b00001100000: begin lvalue_r <= 16'b0000010010110111; rvalue_r <= 16'b0000010011000100;end
            11'b00001100001: begin lvalue_r <= 16'b0000010011000100; rvalue_r <= 16'b0000010011010000;end
            11'b00001100010: begin lvalue_r <= 16'b0000010011010000; rvalue_r <= 16'b0000010011011101;end
            11'b00001100011: begin lvalue_r <= 16'b0000010011011101; rvalue_r <= 16'b0000010011101001;end
            11'b00001100100: begin lvalue_r <= 16'b0000010011101001; rvalue_r <= 16'b0000010011110110;end
            11'b00001100101: begin lvalue_r <= 16'b0000010011110110; rvalue_r <= 16'b0000010100000010;end
            11'b00001100110: begin lvalue_r <= 16'b0000010100000010; rvalue_r <= 16'b0000010100001111;end
            11'b00001100111: begin lvalue_r <= 16'b0000010100001111; rvalue_r <= 16'b0000010100011100;end
            11'b00001101000: begin lvalue_r <= 16'b0000010100011100; rvalue_r <= 16'b0000010100101000;end
            11'b00001101001: begin lvalue_r <= 16'b0000010100101000; rvalue_r <= 16'b0000010100110101;end
            11'b00001101010: begin lvalue_r <= 16'b0000010100110101; rvalue_r <= 16'b0000010101000001;end
            11'b00001101011: begin lvalue_r <= 16'b0000010101000001; rvalue_r <= 16'b0000010101001110;end
            11'b00001101100: begin lvalue_r <= 16'b0000010101001110; rvalue_r <= 16'b0000010101011011;end
            11'b00001101101: begin lvalue_r <= 16'b0000010101011011; rvalue_r <= 16'b0000010101100111;end
            11'b00001101110: begin lvalue_r <= 16'b0000010101100111; rvalue_r <= 16'b0000010101110100;end
            11'b00001101111: begin lvalue_r <= 16'b0000010101110100; rvalue_r <= 16'b0000010110000000;end
            11'b00001110000: begin lvalue_r <= 16'b0000010110000000; rvalue_r <= 16'b0000010110001101;end
            11'b00001110001: begin lvalue_r <= 16'b0000010110001101; rvalue_r <= 16'b0000010110011001;end
            11'b00001110010: begin lvalue_r <= 16'b0000010110011001; rvalue_r <= 16'b0000010110100110;end
            11'b00001110011: begin lvalue_r <= 16'b0000010110100110; rvalue_r <= 16'b0000010110110011;end
            11'b00001110100: begin lvalue_r <= 16'b0000010110110011; rvalue_r <= 16'b0000010110111111;end
            11'b00001110101: begin lvalue_r <= 16'b0000010110111111; rvalue_r <= 16'b0000010111001100;end
            11'b00001110110: begin lvalue_r <= 16'b0000010111001100; rvalue_r <= 16'b0000010111011000;end
            11'b00001110111: begin lvalue_r <= 16'b0000010111011000; rvalue_r <= 16'b0000010111100101;end
            11'b00001111000: begin lvalue_r <= 16'b0000010111100101; rvalue_r <= 16'b0000010111110010;end
            11'b00001111001: begin lvalue_r <= 16'b0000010111110010; rvalue_r <= 16'b0000010111111110;end
            11'b00001111010: begin lvalue_r <= 16'b0000010111111110; rvalue_r <= 16'b0000011000001011;end
            11'b00001111011: begin lvalue_r <= 16'b0000011000001011; rvalue_r <= 16'b0000011000010111;end
            11'b00001111100: begin lvalue_r <= 16'b0000011000010111; rvalue_r <= 16'b0000011000100100;end
            11'b00001111101: begin lvalue_r <= 16'b0000011000100100; rvalue_r <= 16'b0000011000110001;end
            11'b00001111110: begin lvalue_r <= 16'b0000011000110001; rvalue_r <= 16'b0000011000111101;end
            11'b00001111111: begin lvalue_r <= 16'b0000011000111101; rvalue_r <= 16'b0000011001001010;end
            11'b00010000000: begin lvalue_r <= 16'b0000011001001010; rvalue_r <= 16'b0000011001010110;end
            11'b00010000001: begin lvalue_r <= 16'b0000011001010110; rvalue_r <= 16'b0000011001100011;end
            11'b00010000010: begin lvalue_r <= 16'b0000011001100011; rvalue_r <= 16'b0000011001110000;end
            11'b00010000011: begin lvalue_r <= 16'b0000011001110000; rvalue_r <= 16'b0000011001111100;end
            11'b00010000100: begin lvalue_r <= 16'b0000011001111100; rvalue_r <= 16'b0000011010001001;end
            11'b00010000101: begin lvalue_r <= 16'b0000011010001001; rvalue_r <= 16'b0000011010010101;end
            11'b00010000110: begin lvalue_r <= 16'b0000011010010101; rvalue_r <= 16'b0000011010100010;end
            11'b00010000111: begin lvalue_r <= 16'b0000011010100010; rvalue_r <= 16'b0000011010101111;end
            11'b00010001000: begin lvalue_r <= 16'b0000011010101111; rvalue_r <= 16'b0000011010111011;end
            11'b00010001001: begin lvalue_r <= 16'b0000011010111011; rvalue_r <= 16'b0000011011001000;end
            11'b00010001010: begin lvalue_r <= 16'b0000011011001000; rvalue_r <= 16'b0000011011010100;end
            11'b00010001011: begin lvalue_r <= 16'b0000011011010100; rvalue_r <= 16'b0000011011100001;end
            11'b00010001100: begin lvalue_r <= 16'b0000011011100001; rvalue_r <= 16'b0000011011101110;end
            11'b00010001101: begin lvalue_r <= 16'b0000011011101110; rvalue_r <= 16'b0000011011111010;end
            11'b00010001110: begin lvalue_r <= 16'b0000011011111010; rvalue_r <= 16'b0000011100000111;end
            11'b00010001111: begin lvalue_r <= 16'b0000011100000111; rvalue_r <= 16'b0000011100010011;end
            11'b00010010000: begin lvalue_r <= 16'b0000011100010011; rvalue_r <= 16'b0000011100100000;end
            11'b00010010001: begin lvalue_r <= 16'b0000011100100000; rvalue_r <= 16'b0000011100101101;end
            11'b00010010010: begin lvalue_r <= 16'b0000011100101101; rvalue_r <= 16'b0000011100111001;end
            11'b00010010011: begin lvalue_r <= 16'b0000011100111001; rvalue_r <= 16'b0000011101000110;end
            11'b00010010100: begin lvalue_r <= 16'b0000011101000110; rvalue_r <= 16'b0000011101010010;end
            11'b00010010101: begin lvalue_r <= 16'b0000011101010010; rvalue_r <= 16'b0000011101011111;end
            11'b00010010110: begin lvalue_r <= 16'b0000011101011111; rvalue_r <= 16'b0000011101101100;end
            11'b00010010111: begin lvalue_r <= 16'b0000011101101100; rvalue_r <= 16'b0000011101111000;end
            11'b00010011000: begin lvalue_r <= 16'b0000011101111000; rvalue_r <= 16'b0000011110000101;end
            11'b00010011001: begin lvalue_r <= 16'b0000011110000101; rvalue_r <= 16'b0000011110010001;end
            11'b00010011010: begin lvalue_r <= 16'b0000011110010001; rvalue_r <= 16'b0000011110011110;end
            11'b00010011011: begin lvalue_r <= 16'b0000011110011110; rvalue_r <= 16'b0000011110101011;end
            11'b00010011100: begin lvalue_r <= 16'b0000011110101011; rvalue_r <= 16'b0000011110110111;end
            11'b00010011101: begin lvalue_r <= 16'b0000011110110111; rvalue_r <= 16'b0000011111000100;end
            11'b00010011110: begin lvalue_r <= 16'b0000011111000100; rvalue_r <= 16'b0000011111010001;end
            11'b00010011111: begin lvalue_r <= 16'b0000011111010001; rvalue_r <= 16'b0000011111011101;end
            11'b00010100000: begin lvalue_r <= 16'b0000011111011101; rvalue_r <= 16'b0000011111101010;end
            11'b00010100001: begin lvalue_r <= 16'b0000011111101010; rvalue_r <= 16'b0000011111110110;end
            11'b00010100010: begin lvalue_r <= 16'b0000011111110110; rvalue_r <= 16'b0000100000000011;end
            11'b00010100011: begin lvalue_r <= 16'b0000100000000011; rvalue_r <= 16'b0000100000010000;end
            11'b00010100100: begin lvalue_r <= 16'b0000100000010000; rvalue_r <= 16'b0000100000011100;end
            11'b00010100101: begin lvalue_r <= 16'b0000100000011100; rvalue_r <= 16'b0000100000101001;end
            11'b00010100110: begin lvalue_r <= 16'b0000100000101001; rvalue_r <= 16'b0000100000110101;end
            11'b00010100111: begin lvalue_r <= 16'b0000100000110101; rvalue_r <= 16'b0000100001000010;end
            11'b00010101000: begin lvalue_r <= 16'b0000100001000010; rvalue_r <= 16'b0000100001001111;end
            11'b00010101001: begin lvalue_r <= 16'b0000100001001111; rvalue_r <= 16'b0000100001011011;end
            11'b00010101010: begin lvalue_r <= 16'b0000100001011011; rvalue_r <= 16'b0000100001101000;end
            11'b00010101011: begin lvalue_r <= 16'b0000100001101000; rvalue_r <= 16'b0000100001110101;end
            11'b00010101100: begin lvalue_r <= 16'b0000100001110101; rvalue_r <= 16'b0000100010000001;end
            11'b00010101101: begin lvalue_r <= 16'b0000100010000001; rvalue_r <= 16'b0000100010001110;end
            11'b00010101110: begin lvalue_r <= 16'b0000100010001110; rvalue_r <= 16'b0000100010011010;end
            11'b00010101111: begin lvalue_r <= 16'b0000100010011010; rvalue_r <= 16'b0000100010100111;end
            11'b00010110000: begin lvalue_r <= 16'b0000100010100111; rvalue_r <= 16'b0000100010110100;end
            11'b00010110001: begin lvalue_r <= 16'b0000100010110100; rvalue_r <= 16'b0000100011000000;end
            11'b00010110010: begin lvalue_r <= 16'b0000100011000000; rvalue_r <= 16'b0000100011001101;end
            11'b00010110011: begin lvalue_r <= 16'b0000100011001101; rvalue_r <= 16'b0000100011011010;end
            11'b00010110100: begin lvalue_r <= 16'b0000100011011010; rvalue_r <= 16'b0000100011100110;end
            11'b00010110101: begin lvalue_r <= 16'b0000100011100110; rvalue_r <= 16'b0000100011110011;end
            11'b00010110110: begin lvalue_r <= 16'b0000100011110011; rvalue_r <= 16'b0000100011111111;end
            11'b00010110111: begin lvalue_r <= 16'b0000100011111111; rvalue_r <= 16'b0000100100001100;end
            11'b00010111000: begin lvalue_r <= 16'b0000100100001100; rvalue_r <= 16'b0000100100011001;end
            11'b00010111001: begin lvalue_r <= 16'b0000100100011001; rvalue_r <= 16'b0000100100100101;end
            11'b00010111010: begin lvalue_r <= 16'b0000100100100101; rvalue_r <= 16'b0000100100110010;end
            11'b00010111011: begin lvalue_r <= 16'b0000100100110010; rvalue_r <= 16'b0000100100111111;end
            11'b00010111100: begin lvalue_r <= 16'b0000100100111111; rvalue_r <= 16'b0000100101001011;end
            11'b00010111101: begin lvalue_r <= 16'b0000100101001011; rvalue_r <= 16'b0000100101011000;end
            11'b00010111110: begin lvalue_r <= 16'b0000100101011000; rvalue_r <= 16'b0000100101100100;end
            11'b00010111111: begin lvalue_r <= 16'b0000100101100100; rvalue_r <= 16'b0000100101110001;end
            11'b00011000000: begin lvalue_r <= 16'b0000100101110001; rvalue_r <= 16'b0000100101111110;end
            11'b00011000001: begin lvalue_r <= 16'b0000100101111110; rvalue_r <= 16'b0000100110001010;end
            11'b00011000010: begin lvalue_r <= 16'b0000100110001010; rvalue_r <= 16'b0000100110010111;end
            11'b00011000011: begin lvalue_r <= 16'b0000100110010111; rvalue_r <= 16'b0000100110100100;end
            11'b00011000100: begin lvalue_r <= 16'b0000100110100100; rvalue_r <= 16'b0000100110110000;end
            11'b00011000101: begin lvalue_r <= 16'b0000100110110000; rvalue_r <= 16'b0000100110111101;end
            11'b00011000110: begin lvalue_r <= 16'b0000100110111101; rvalue_r <= 16'b0000100111001010;end
            11'b00011000111: begin lvalue_r <= 16'b0000100111001010; rvalue_r <= 16'b0000100111010110;end
            11'b00011001000: begin lvalue_r <= 16'b0000100111010110; rvalue_r <= 16'b0000100111100011;end
            11'b00011001001: begin lvalue_r <= 16'b0000100111100011; rvalue_r <= 16'b0000100111101111;end
            11'b00011001010: begin lvalue_r <= 16'b0000100111101111; rvalue_r <= 16'b0000100111111100;end
            11'b00011001011: begin lvalue_r <= 16'b0000100111111100; rvalue_r <= 16'b0000101000001001;end
            11'b00011001100: begin lvalue_r <= 16'b0000101000001001; rvalue_r <= 16'b0000101000010101;end
            11'b00011001101: begin lvalue_r <= 16'b0000101000010101; rvalue_r <= 16'b0000101000100010;end
            11'b00011001110: begin lvalue_r <= 16'b0000101000100010; rvalue_r <= 16'b0000101000101111;end
            11'b00011001111: begin lvalue_r <= 16'b0000101000101111; rvalue_r <= 16'b0000101000111011;end
            11'b00011010000: begin lvalue_r <= 16'b0000101000111011; rvalue_r <= 16'b0000101001001000;end
            11'b00011010001: begin lvalue_r <= 16'b0000101001001000; rvalue_r <= 16'b0000101001010101;end
            11'b00011010010: begin lvalue_r <= 16'b0000101001010101; rvalue_r <= 16'b0000101001100001;end
            11'b00011010011: begin lvalue_r <= 16'b0000101001100001; rvalue_r <= 16'b0000101001101110;end
            11'b00011010100: begin lvalue_r <= 16'b0000101001101110; rvalue_r <= 16'b0000101001111011;end
            11'b00011010101: begin lvalue_r <= 16'b0000101001111011; rvalue_r <= 16'b0000101010000111;end
            11'b00011010110: begin lvalue_r <= 16'b0000101010000111; rvalue_r <= 16'b0000101010010100;end
            11'b00011010111: begin lvalue_r <= 16'b0000101010010100; rvalue_r <= 16'b0000101010100001;end
            11'b00011011000: begin lvalue_r <= 16'b0000101010100001; rvalue_r <= 16'b0000101010101101;end
            11'b00011011001: begin lvalue_r <= 16'b0000101010101101; rvalue_r <= 16'b0000101010111010;end
            11'b00011011010: begin lvalue_r <= 16'b0000101010111010; rvalue_r <= 16'b0000101011000111;end
            11'b00011011011: begin lvalue_r <= 16'b0000101011000111; rvalue_r <= 16'b0000101011010011;end
            11'b00011011100: begin lvalue_r <= 16'b0000101011010011; rvalue_r <= 16'b0000101011100000;end
            11'b00011011101: begin lvalue_r <= 16'b0000101011100000; rvalue_r <= 16'b0000101011101100;end
            11'b00011011110: begin lvalue_r <= 16'b0000101011101100; rvalue_r <= 16'b0000101011111001;end
            11'b00011011111: begin lvalue_r <= 16'b0000101011111001; rvalue_r <= 16'b0000101100000110;end
            11'b00011100000: begin lvalue_r <= 16'b0000101100000110; rvalue_r <= 16'b0000101100010010;end
            11'b00011100001: begin lvalue_r <= 16'b0000101100010010; rvalue_r <= 16'b0000101100011111;end
            11'b00011100010: begin lvalue_r <= 16'b0000101100011111; rvalue_r <= 16'b0000101100101100;end
            11'b00011100011: begin lvalue_r <= 16'b0000101100101100; rvalue_r <= 16'b0000101100111000;end
            11'b00011100100: begin lvalue_r <= 16'b0000101100111000; rvalue_r <= 16'b0000101101000101;end
            11'b00011100101: begin lvalue_r <= 16'b0000101101000101; rvalue_r <= 16'b0000101101010010;end
            11'b00011100110: begin lvalue_r <= 16'b0000101101010010; rvalue_r <= 16'b0000101101011110;end
            11'b00011100111: begin lvalue_r <= 16'b0000101101011110; rvalue_r <= 16'b0000101101101011;end
            11'b00011101000: begin lvalue_r <= 16'b0000101101101011; rvalue_r <= 16'b0000101101111000;end
            11'b00011101001: begin lvalue_r <= 16'b0000101101111000; rvalue_r <= 16'b0000101110000100;end
            11'b00011101010: begin lvalue_r <= 16'b0000101110000100; rvalue_r <= 16'b0000101110010001;end
            11'b00011101011: begin lvalue_r <= 16'b0000101110010001; rvalue_r <= 16'b0000101110011110;end
            11'b00011101100: begin lvalue_r <= 16'b0000101110011110; rvalue_r <= 16'b0000101110101010;end
            11'b00011101101: begin lvalue_r <= 16'b0000101110101010; rvalue_r <= 16'b0000101110110111;end
            11'b00011101110: begin lvalue_r <= 16'b0000101110110111; rvalue_r <= 16'b0000101111000100;end
            11'b00011101111: begin lvalue_r <= 16'b0000101111000100; rvalue_r <= 16'b0000101111010000;end
            11'b00011110000: begin lvalue_r <= 16'b0000101111010000; rvalue_r <= 16'b0000101111011101;end
            11'b00011110001: begin lvalue_r <= 16'b0000101111011101; rvalue_r <= 16'b0000101111101010;end
            11'b00011110010: begin lvalue_r <= 16'b0000101111101010; rvalue_r <= 16'b0000101111110110;end
            11'b00011110011: begin lvalue_r <= 16'b0000101111110110; rvalue_r <= 16'b0000110000000011;end
            11'b00011110100: begin lvalue_r <= 16'b0000110000000011; rvalue_r <= 16'b0000110000010000;end
            11'b00011110101: begin lvalue_r <= 16'b0000110000010000; rvalue_r <= 16'b0000110000011101;end
            11'b00011110110: begin lvalue_r <= 16'b0000110000011101; rvalue_r <= 16'b0000110000101001;end
            11'b00011110111: begin lvalue_r <= 16'b0000110000101001; rvalue_r <= 16'b0000110000110110;end
            11'b00011111000: begin lvalue_r <= 16'b0000110000110110; rvalue_r <= 16'b0000110001000011;end
            11'b00011111001: begin lvalue_r <= 16'b0000110001000011; rvalue_r <= 16'b0000110001001111;end
            11'b00011111010: begin lvalue_r <= 16'b0000110001001111; rvalue_r <= 16'b0000110001011100;end
            11'b00011111011: begin lvalue_r <= 16'b0000110001011100; rvalue_r <= 16'b0000110001101001;end
            11'b00011111100: begin lvalue_r <= 16'b0000110001101001; rvalue_r <= 16'b0000110001110101;end
            11'b00011111101: begin lvalue_r <= 16'b0000110001110101; rvalue_r <= 16'b0000110010000010;end
            11'b00011111110: begin lvalue_r <= 16'b0000110010000010; rvalue_r <= 16'b0000110010001111;end
            11'b00011111111: begin lvalue_r <= 16'b0000110010001111; rvalue_r <= 16'b0000110010011011;end
            11'b00100000000: begin lvalue_r <= 16'b0000110010011011; rvalue_r <= 16'b0000110010101000;end
            11'b00100000001: begin lvalue_r <= 16'b0000110010101000; rvalue_r <= 16'b0000110010110101;end
            11'b00100000010: begin lvalue_r <= 16'b0000110010110101; rvalue_r <= 16'b0000110011000001;end
            11'b00100000011: begin lvalue_r <= 16'b0000110011000001; rvalue_r <= 16'b0000110011001110;end
            11'b00100000100: begin lvalue_r <= 16'b0000110011001110; rvalue_r <= 16'b0000110011011011;end
            11'b00100000101: begin lvalue_r <= 16'b0000110011011011; rvalue_r <= 16'b0000110011101000;end
            11'b00100000110: begin lvalue_r <= 16'b0000110011101000; rvalue_r <= 16'b0000110011110100;end
            11'b00100000111: begin lvalue_r <= 16'b0000110011110100; rvalue_r <= 16'b0000110100000001;end
            11'b00100001000: begin lvalue_r <= 16'b0000110100000001; rvalue_r <= 16'b0000110100001110;end
            11'b00100001001: begin lvalue_r <= 16'b0000110100001110; rvalue_r <= 16'b0000110100011010;end
            11'b00100001010: begin lvalue_r <= 16'b0000110100011010; rvalue_r <= 16'b0000110100100111;end
            11'b00100001011: begin lvalue_r <= 16'b0000110100100111; rvalue_r <= 16'b0000110100110100;end
            11'b00100001100: begin lvalue_r <= 16'b0000110100110100; rvalue_r <= 16'b0000110101000000;end
            11'b00100001101: begin lvalue_r <= 16'b0000110101000000; rvalue_r <= 16'b0000110101001101;end
            11'b00100001110: begin lvalue_r <= 16'b0000110101001101; rvalue_r <= 16'b0000110101011010;end
            11'b00100001111: begin lvalue_r <= 16'b0000110101011010; rvalue_r <= 16'b0000110101100111;end
            11'b00100010000: begin lvalue_r <= 16'b0000110101100111; rvalue_r <= 16'b0000110101110011;end
            11'b00100010001: begin lvalue_r <= 16'b0000110101110011; rvalue_r <= 16'b0000110110000000;end
            11'b00100010010: begin lvalue_r <= 16'b0000110110000000; rvalue_r <= 16'b0000110110001101;end
            11'b00100010011: begin lvalue_r <= 16'b0000110110001101; rvalue_r <= 16'b0000110110011001;end
            11'b00100010100: begin lvalue_r <= 16'b0000110110011001; rvalue_r <= 16'b0000110110100110;end
            11'b00100010101: begin lvalue_r <= 16'b0000110110100110; rvalue_r <= 16'b0000110110110011;end
            11'b00100010110: begin lvalue_r <= 16'b0000110110110011; rvalue_r <= 16'b0000110110111111;end
            11'b00100010111: begin lvalue_r <= 16'b0000110110111111; rvalue_r <= 16'b0000110111001100;end
            11'b00100011000: begin lvalue_r <= 16'b0000110111001100; rvalue_r <= 16'b0000110111011001;end
            11'b00100011001: begin lvalue_r <= 16'b0000110111011001; rvalue_r <= 16'b0000110111100110;end
            11'b00100011010: begin lvalue_r <= 16'b0000110111100110; rvalue_r <= 16'b0000110111110010;end
            11'b00100011011: begin lvalue_r <= 16'b0000110111110010; rvalue_r <= 16'b0000110111111111;end
            11'b00100011100: begin lvalue_r <= 16'b0000110111111111; rvalue_r <= 16'b0000111000001100;end
            11'b00100011101: begin lvalue_r <= 16'b0000111000001100; rvalue_r <= 16'b0000111000011000;end
            11'b00100011110: begin lvalue_r <= 16'b0000111000011000; rvalue_r <= 16'b0000111000100101;end
            11'b00100011111: begin lvalue_r <= 16'b0000111000100101; rvalue_r <= 16'b0000111000110010;end
            11'b00100100000: begin lvalue_r <= 16'b0000111000110010; rvalue_r <= 16'b0000111000111111;end
            11'b00100100001: begin lvalue_r <= 16'b0000111000111111; rvalue_r <= 16'b0000111001001011;end
            11'b00100100010: begin lvalue_r <= 16'b0000111001001011; rvalue_r <= 16'b0000111001011000;end
            11'b00100100011: begin lvalue_r <= 16'b0000111001011000; rvalue_r <= 16'b0000111001100101;end
            11'b00100100100: begin lvalue_r <= 16'b0000111001100101; rvalue_r <= 16'b0000111001110010;end
            11'b00100100101: begin lvalue_r <= 16'b0000111001110010; rvalue_r <= 16'b0000111001111110;end
            11'b00100100110: begin lvalue_r <= 16'b0000111001111110; rvalue_r <= 16'b0000111010001011;end
            11'b00100100111: begin lvalue_r <= 16'b0000111010001011; rvalue_r <= 16'b0000111010011000;end
            11'b00100101000: begin lvalue_r <= 16'b0000111010011000; rvalue_r <= 16'b0000111010100100;end
            11'b00100101001: begin lvalue_r <= 16'b0000111010100100; rvalue_r <= 16'b0000111010110001;end
            11'b00100101010: begin lvalue_r <= 16'b0000111010110001; rvalue_r <= 16'b0000111010111110;end
            11'b00100101011: begin lvalue_r <= 16'b0000111010111110; rvalue_r <= 16'b0000111011001011;end
            11'b00100101100: begin lvalue_r <= 16'b0000111011001011; rvalue_r <= 16'b0000111011010111;end
            11'b00100101101: begin lvalue_r <= 16'b0000111011010111; rvalue_r <= 16'b0000111011100100;end
            11'b00100101110: begin lvalue_r <= 16'b0000111011100100; rvalue_r <= 16'b0000111011110001;end
            11'b00100101111: begin lvalue_r <= 16'b0000111011110001; rvalue_r <= 16'b0000111011111110;end
            11'b00100110000: begin lvalue_r <= 16'b0000111011111110; rvalue_r <= 16'b0000111100001010;end
            11'b00100110001: begin lvalue_r <= 16'b0000111100001010; rvalue_r <= 16'b0000111100010111;end
            11'b00100110010: begin lvalue_r <= 16'b0000111100010111; rvalue_r <= 16'b0000111100100100;end
            11'b00100110011: begin lvalue_r <= 16'b0000111100100100; rvalue_r <= 16'b0000111100110001;end
            11'b00100110100: begin lvalue_r <= 16'b0000111100110001; rvalue_r <= 16'b0000111100111101;end
            11'b00100110101: begin lvalue_r <= 16'b0000111100111101; rvalue_r <= 16'b0000111101001010;end
            11'b00100110110: begin lvalue_r <= 16'b0000111101001010; rvalue_r <= 16'b0000111101010111;end
            11'b00100110111: begin lvalue_r <= 16'b0000111101010111; rvalue_r <= 16'b0000111101100100;end
            11'b00100111000: begin lvalue_r <= 16'b0000111101100100; rvalue_r <= 16'b0000111101110000;end
            11'b00100111001: begin lvalue_r <= 16'b0000111101110000; rvalue_r <= 16'b0000111101111101;end
            11'b00100111010: begin lvalue_r <= 16'b0000111101111101; rvalue_r <= 16'b0000111110001010;end
            11'b00100111011: begin lvalue_r <= 16'b0000111110001010; rvalue_r <= 16'b0000111110010111;end
            11'b00100111100: begin lvalue_r <= 16'b0000111110010111; rvalue_r <= 16'b0000111110100011;end
            11'b00100111101: begin lvalue_r <= 16'b0000111110100011; rvalue_r <= 16'b0000111110110000;end
            11'b00100111110: begin lvalue_r <= 16'b0000111110110000; rvalue_r <= 16'b0000111110111101;end
            11'b00100111111: begin lvalue_r <= 16'b0000111110111101; rvalue_r <= 16'b0000111111001010;end
            11'b00101000000: begin lvalue_r <= 16'b0000111111001010; rvalue_r <= 16'b0000111111010110;end
            11'b00101000001: begin lvalue_r <= 16'b0000111111010110; rvalue_r <= 16'b0000111111100011;end
            11'b00101000010: begin lvalue_r <= 16'b0000111111100011; rvalue_r <= 16'b0000111111110000;end
            11'b00101000011: begin lvalue_r <= 16'b0000111111110000; rvalue_r <= 16'b0000111111111101;end
            11'b00101000100: begin lvalue_r <= 16'b0000111111111101; rvalue_r <= 16'b0001000000001001;end
            11'b00101000101: begin lvalue_r <= 16'b0001000000001001; rvalue_r <= 16'b0001000000010110;end
            11'b00101000110: begin lvalue_r <= 16'b0001000000010110; rvalue_r <= 16'b0001000000100011;end
            11'b00101000111: begin lvalue_r <= 16'b0001000000100011; rvalue_r <= 16'b0001000000110000;end
            11'b00101001000: begin lvalue_r <= 16'b0001000000110000; rvalue_r <= 16'b0001000000111100;end
            11'b00101001001: begin lvalue_r <= 16'b0001000000111100; rvalue_r <= 16'b0001000001001001;end
            11'b00101001010: begin lvalue_r <= 16'b0001000001001001; rvalue_r <= 16'b0001000001010110;end
            11'b00101001011: begin lvalue_r <= 16'b0001000001010110; rvalue_r <= 16'b0001000001100011;end
            11'b00101001100: begin lvalue_r <= 16'b0001000001100011; rvalue_r <= 16'b0001000001101111;end
            11'b00101001101: begin lvalue_r <= 16'b0001000001101111; rvalue_r <= 16'b0001000001111100;end
            11'b00101001110: begin lvalue_r <= 16'b0001000001111100; rvalue_r <= 16'b0001000010001001;end
            11'b00101001111: begin lvalue_r <= 16'b0001000010001001; rvalue_r <= 16'b0001000010010110;end
            11'b00101010000: begin lvalue_r <= 16'b0001000010010110; rvalue_r <= 16'b0001000010100011;end
            11'b00101010001: begin lvalue_r <= 16'b0001000010100011; rvalue_r <= 16'b0001000010101111;end
            11'b00101010010: begin lvalue_r <= 16'b0001000010101111; rvalue_r <= 16'b0001000010111100;end
            11'b00101010011: begin lvalue_r <= 16'b0001000010111100; rvalue_r <= 16'b0001000011001001;end
            11'b00101010100: begin lvalue_r <= 16'b0001000011001001; rvalue_r <= 16'b0001000011010110;end
            11'b00101010101: begin lvalue_r <= 16'b0001000011010110; rvalue_r <= 16'b0001000011100011;end
            11'b00101010110: begin lvalue_r <= 16'b0001000011100011; rvalue_r <= 16'b0001000011101111;end
            11'b00101010111: begin lvalue_r <= 16'b0001000011101111; rvalue_r <= 16'b0001000011111100;end
            11'b00101011000: begin lvalue_r <= 16'b0001000011111100; rvalue_r <= 16'b0001000100001001;end
            11'b00101011001: begin lvalue_r <= 16'b0001000100001001; rvalue_r <= 16'b0001000100010110;end
            11'b00101011010: begin lvalue_r <= 16'b0001000100010110; rvalue_r <= 16'b0001000100100010;end
            11'b00101011011: begin lvalue_r <= 16'b0001000100100010; rvalue_r <= 16'b0001000100101111;end
            11'b00101011100: begin lvalue_r <= 16'b0001000100101111; rvalue_r <= 16'b0001000100111100;end
            11'b00101011101: begin lvalue_r <= 16'b0001000100111100; rvalue_r <= 16'b0001000101001001;end
            11'b00101011110: begin lvalue_r <= 16'b0001000101001001; rvalue_r <= 16'b0001000101010110;end
            11'b00101011111: begin lvalue_r <= 16'b0001000101010110; rvalue_r <= 16'b0001000101100010;end
            11'b00101100000: begin lvalue_r <= 16'b0001000101100010; rvalue_r <= 16'b0001000101101111;end
            11'b00101100001: begin lvalue_r <= 16'b0001000101101111; rvalue_r <= 16'b0001000101111100;end
            11'b00101100010: begin lvalue_r <= 16'b0001000101111100; rvalue_r <= 16'b0001000110001001;end
            11'b00101100011: begin lvalue_r <= 16'b0001000110001001; rvalue_r <= 16'b0001000110010110;end
            11'b00101100100: begin lvalue_r <= 16'b0001000110010110; rvalue_r <= 16'b0001000110100010;end
            11'b00101100101: begin lvalue_r <= 16'b0001000110100010; rvalue_r <= 16'b0001000110101111;end
            11'b00101100110: begin lvalue_r <= 16'b0001000110101111; rvalue_r <= 16'b0001000110111100;end
            11'b00101100111: begin lvalue_r <= 16'b0001000110111100; rvalue_r <= 16'b0001000111001001;end
            11'b00101101000: begin lvalue_r <= 16'b0001000111001001; rvalue_r <= 16'b0001000111010110;end
            11'b00101101001: begin lvalue_r <= 16'b0001000111010110; rvalue_r <= 16'b0001000111100010;end
            11'b00101101010: begin lvalue_r <= 16'b0001000111100010; rvalue_r <= 16'b0001000111101111;end
            11'b00101101011: begin lvalue_r <= 16'b0001000111101111; rvalue_r <= 16'b0001000111111100;end
            11'b00101101100: begin lvalue_r <= 16'b0001000111111100; rvalue_r <= 16'b0001001000001001;end
            11'b00101101101: begin lvalue_r <= 16'b0001001000001001; rvalue_r <= 16'b0001001000010110;end
            11'b00101101110: begin lvalue_r <= 16'b0001001000010110; rvalue_r <= 16'b0001001000100011;end
            11'b00101101111: begin lvalue_r <= 16'b0001001000100011; rvalue_r <= 16'b0001001000101111;end
            11'b00101110000: begin lvalue_r <= 16'b0001001000101111; rvalue_r <= 16'b0001001000111100;end
            11'b00101110001: begin lvalue_r <= 16'b0001001000111100; rvalue_r <= 16'b0001001001001001;end
            11'b00101110010: begin lvalue_r <= 16'b0001001001001001; rvalue_r <= 16'b0001001001010110;end
            11'b00101110011: begin lvalue_r <= 16'b0001001001010110; rvalue_r <= 16'b0001001001100011;end
            11'b00101110100: begin lvalue_r <= 16'b0001001001100011; rvalue_r <= 16'b0001001001101111;end
            11'b00101110101: begin lvalue_r <= 16'b0001001001101111; rvalue_r <= 16'b0001001001111100;end
            11'b00101110110: begin lvalue_r <= 16'b0001001001111100; rvalue_r <= 16'b0001001010001001;end
            11'b00101110111: begin lvalue_r <= 16'b0001001010001001; rvalue_r <= 16'b0001001010010110;end
            11'b00101111000: begin lvalue_r <= 16'b0001001010010110; rvalue_r <= 16'b0001001010100011;end
            11'b00101111001: begin lvalue_r <= 16'b0001001010100011; rvalue_r <= 16'b0001001010110000;end
            11'b00101111010: begin lvalue_r <= 16'b0001001010110000; rvalue_r <= 16'b0001001010111100;end
            11'b00101111011: begin lvalue_r <= 16'b0001001010111100; rvalue_r <= 16'b0001001011001001;end
            11'b00101111100: begin lvalue_r <= 16'b0001001011001001; rvalue_r <= 16'b0001001011010110;end
            11'b00101111101: begin lvalue_r <= 16'b0001001011010110; rvalue_r <= 16'b0001001011100011;end
            11'b00101111110: begin lvalue_r <= 16'b0001001011100011; rvalue_r <= 16'b0001001011110000;end
            11'b00101111111: begin lvalue_r <= 16'b0001001011110000; rvalue_r <= 16'b0001001011111101;end
            11'b00110000000: begin lvalue_r <= 16'b0001001011111101; rvalue_r <= 16'b0001001100001010;end
            11'b00110000001: begin lvalue_r <= 16'b0001001100001010; rvalue_r <= 16'b0001001100010110;end
            11'b00110000010: begin lvalue_r <= 16'b0001001100010110; rvalue_r <= 16'b0001001100100011;end
            11'b00110000011: begin lvalue_r <= 16'b0001001100100011; rvalue_r <= 16'b0001001100110000;end
            11'b00110000100: begin lvalue_r <= 16'b0001001100110000; rvalue_r <= 16'b0001001100111101;end
            11'b00110000101: begin lvalue_r <= 16'b0001001100111101; rvalue_r <= 16'b0001001101001010;end
            11'b00110000110: begin lvalue_r <= 16'b0001001101001010; rvalue_r <= 16'b0001001101010111;end
            11'b00110000111: begin lvalue_r <= 16'b0001001101010111; rvalue_r <= 16'b0001001101100011;end
            11'b00110001000: begin lvalue_r <= 16'b0001001101100011; rvalue_r <= 16'b0001001101110000;end
            11'b00110001001: begin lvalue_r <= 16'b0001001101110000; rvalue_r <= 16'b0001001101111101;end
            11'b00110001010: begin lvalue_r <= 16'b0001001101111101; rvalue_r <= 16'b0001001110001010;end
            11'b00110001011: begin lvalue_r <= 16'b0001001110001010; rvalue_r <= 16'b0001001110010111;end
            11'b00110001100: begin lvalue_r <= 16'b0001001110010111; rvalue_r <= 16'b0001001110100100;end
            11'b00110001101: begin lvalue_r <= 16'b0001001110100100; rvalue_r <= 16'b0001001110110001;end
            11'b00110001110: begin lvalue_r <= 16'b0001001110110001; rvalue_r <= 16'b0001001110111101;end
            11'b00110001111: begin lvalue_r <= 16'b0001001110111101; rvalue_r <= 16'b0001001111001010;end
            11'b00110010000: begin lvalue_r <= 16'b0001001111001010; rvalue_r <= 16'b0001001111010111;end
            11'b00110010001: begin lvalue_r <= 16'b0001001111010111; rvalue_r <= 16'b0001001111100100;end
            11'b00110010010: begin lvalue_r <= 16'b0001001111100100; rvalue_r <= 16'b0001001111110001;end
            11'b00110010011: begin lvalue_r <= 16'b0001001111110001; rvalue_r <= 16'b0001001111111110;end
            11'b00110010100: begin lvalue_r <= 16'b0001001111111110; rvalue_r <= 16'b0001010000001011;end
            11'b00110010101: begin lvalue_r <= 16'b0001010000001011; rvalue_r <= 16'b0001010000011000;end
            11'b00110010110: begin lvalue_r <= 16'b0001010000011000; rvalue_r <= 16'b0001010000100100;end
            11'b00110010111: begin lvalue_r <= 16'b0001010000100100; rvalue_r <= 16'b0001010000110001;end
            11'b00110011000: begin lvalue_r <= 16'b0001010000110001; rvalue_r <= 16'b0001010000111110;end
            11'b00110011001: begin lvalue_r <= 16'b0001010000111110; rvalue_r <= 16'b0001010001001011;end
            11'b00110011010: begin lvalue_r <= 16'b0001010001001011; rvalue_r <= 16'b0001010001011000;end
            11'b00110011011: begin lvalue_r <= 16'b0001010001011000; rvalue_r <= 16'b0001010001100101;end
            11'b00110011100: begin lvalue_r <= 16'b0001010001100101; rvalue_r <= 16'b0001010001110010;end
            11'b00110011101: begin lvalue_r <= 16'b0001010001110010; rvalue_r <= 16'b0001010001111111;end
            11'b00110011110: begin lvalue_r <= 16'b0001010001111111; rvalue_r <= 16'b0001010010001100;end
            11'b00110011111: begin lvalue_r <= 16'b0001010010001100; rvalue_r <= 16'b0001010010011000;end
            11'b00110100000: begin lvalue_r <= 16'b0001010010011000; rvalue_r <= 16'b0001010010100101;end
            11'b00110100001: begin lvalue_r <= 16'b0001010010100101; rvalue_r <= 16'b0001010010110010;end
            11'b00110100010: begin lvalue_r <= 16'b0001010010110010; rvalue_r <= 16'b0001010010111111;end
            11'b00110100011: begin lvalue_r <= 16'b0001010010111111; rvalue_r <= 16'b0001010011001100;end
            11'b00110100100: begin lvalue_r <= 16'b0001010011001100; rvalue_r <= 16'b0001010011011001;end
            11'b00110100101: begin lvalue_r <= 16'b0001010011011001; rvalue_r <= 16'b0001010011100110;end
            11'b00110100110: begin lvalue_r <= 16'b0001010011100110; rvalue_r <= 16'b0001010011110011;end
            11'b00110100111: begin lvalue_r <= 16'b0001010011110011; rvalue_r <= 16'b0001010100000000;end
            11'b00110101000: begin lvalue_r <= 16'b0001010100000000; rvalue_r <= 16'b0001010100001101;end
            11'b00110101001: begin lvalue_r <= 16'b0001010100001101; rvalue_r <= 16'b0001010100011001;end
            11'b00110101010: begin lvalue_r <= 16'b0001010100011001; rvalue_r <= 16'b0001010100100110;end
            11'b00110101011: begin lvalue_r <= 16'b0001010100100110; rvalue_r <= 16'b0001010100110011;end
            11'b00110101100: begin lvalue_r <= 16'b0001010100110011; rvalue_r <= 16'b0001010101000000;end
            11'b00110101101: begin lvalue_r <= 16'b0001010101000000; rvalue_r <= 16'b0001010101001101;end
            11'b00110101110: begin lvalue_r <= 16'b0001010101001101; rvalue_r <= 16'b0001010101011010;end
            11'b00110101111: begin lvalue_r <= 16'b0001010101011010; rvalue_r <= 16'b0001010101100111;end
            11'b00110110000: begin lvalue_r <= 16'b0001010101100111; rvalue_r <= 16'b0001010101110100;end
            11'b00110110001: begin lvalue_r <= 16'b0001010101110100; rvalue_r <= 16'b0001010110000001;end
            11'b00110110010: begin lvalue_r <= 16'b0001010110000001; rvalue_r <= 16'b0001010110001110;end
            11'b00110110011: begin lvalue_r <= 16'b0001010110001110; rvalue_r <= 16'b0001010110011011;end
            11'b00110110100: begin lvalue_r <= 16'b0001010110011011; rvalue_r <= 16'b0001010110100111;end
            11'b00110110101: begin lvalue_r <= 16'b0001010110100111; rvalue_r <= 16'b0001010110110100;end
            11'b00110110110: begin lvalue_r <= 16'b0001010110110100; rvalue_r <= 16'b0001010111000001;end
            11'b00110110111: begin lvalue_r <= 16'b0001010111000001; rvalue_r <= 16'b0001010111001110;end
            11'b00110111000: begin lvalue_r <= 16'b0001010111001110; rvalue_r <= 16'b0001010111011011;end
            11'b00110111001: begin lvalue_r <= 16'b0001010111011011; rvalue_r <= 16'b0001010111101000;end
            11'b00110111010: begin lvalue_r <= 16'b0001010111101000; rvalue_r <= 16'b0001010111110101;end
            11'b00110111011: begin lvalue_r <= 16'b0001010111110101; rvalue_r <= 16'b0001011000000010;end
            11'b00110111100: begin lvalue_r <= 16'b0001011000000010; rvalue_r <= 16'b0001011000001111;end
            11'b00110111101: begin lvalue_r <= 16'b0001011000001111; rvalue_r <= 16'b0001011000011100;end
            11'b00110111110: begin lvalue_r <= 16'b0001011000011100; rvalue_r <= 16'b0001011000101001;end
            11'b00110111111: begin lvalue_r <= 16'b0001011000101001; rvalue_r <= 16'b0001011000110110;end
            11'b00111000000: begin lvalue_r <= 16'b0001011000110110; rvalue_r <= 16'b0001011001000011;end
            11'b00111000001: begin lvalue_r <= 16'b0001011001000011; rvalue_r <= 16'b0001011001010000;end
            11'b00111000010: begin lvalue_r <= 16'b0001011001010000; rvalue_r <= 16'b0001011001011101;end
            11'b00111000011: begin lvalue_r <= 16'b0001011001011101; rvalue_r <= 16'b0001011001101010;end
            11'b00111000100: begin lvalue_r <= 16'b0001011001101010; rvalue_r <= 16'b0001011001110111;end
            11'b00111000101: begin lvalue_r <= 16'b0001011001110111; rvalue_r <= 16'b0001011010000011;end
            11'b00111000110: begin lvalue_r <= 16'b0001011010000011; rvalue_r <= 16'b0001011010010000;end
            11'b00111000111: begin lvalue_r <= 16'b0001011010010000; rvalue_r <= 16'b0001011010011101;end
            11'b00111001000: begin lvalue_r <= 16'b0001011010011101; rvalue_r <= 16'b0001011010101010;end
            11'b00111001001: begin lvalue_r <= 16'b0001011010101010; rvalue_r <= 16'b0001011010110111;end
            11'b00111001010: begin lvalue_r <= 16'b0001011010110111; rvalue_r <= 16'b0001011011000100;end
            11'b00111001011: begin lvalue_r <= 16'b0001011011000100; rvalue_r <= 16'b0001011011010001;end
            11'b00111001100: begin lvalue_r <= 16'b0001011011010001; rvalue_r <= 16'b0001011011011110;end
            11'b00111001101: begin lvalue_r <= 16'b0001011011011110; rvalue_r <= 16'b0001011011101011;end
            11'b00111001110: begin lvalue_r <= 16'b0001011011101011; rvalue_r <= 16'b0001011011111000;end
            11'b00111001111: begin lvalue_r <= 16'b0001011011111000; rvalue_r <= 16'b0001011100000101;end
            11'b00111010000: begin lvalue_r <= 16'b0001011100000101; rvalue_r <= 16'b0001011100010010;end
            11'b00111010001: begin lvalue_r <= 16'b0001011100010010; rvalue_r <= 16'b0001011100011111;end
            11'b00111010010: begin lvalue_r <= 16'b0001011100011111; rvalue_r <= 16'b0001011100101100;end
            11'b00111010011: begin lvalue_r <= 16'b0001011100101100; rvalue_r <= 16'b0001011100111001;end
            11'b00111010100: begin lvalue_r <= 16'b0001011100111001; rvalue_r <= 16'b0001011101000110;end
            11'b00111010101: begin lvalue_r <= 16'b0001011101000110; rvalue_r <= 16'b0001011101010011;end
            11'b00111010110: begin lvalue_r <= 16'b0001011101010011; rvalue_r <= 16'b0001011101100000;end
            11'b00111010111: begin lvalue_r <= 16'b0001011101100000; rvalue_r <= 16'b0001011101101101;end
            11'b00111011000: begin lvalue_r <= 16'b0001011101101101; rvalue_r <= 16'b0001011101111010;end
            11'b00111011001: begin lvalue_r <= 16'b0001011101111010; rvalue_r <= 16'b0001011110000111;end
            11'b00111011010: begin lvalue_r <= 16'b0001011110000111; rvalue_r <= 16'b0001011110010100;end
            11'b00111011011: begin lvalue_r <= 16'b0001011110010100; rvalue_r <= 16'b0001011110100001;end
            11'b00111011100: begin lvalue_r <= 16'b0001011110100001; rvalue_r <= 16'b0001011110101110;end
            11'b00111011101: begin lvalue_r <= 16'b0001011110101110; rvalue_r <= 16'b0001011110111011;end
            11'b00111011110: begin lvalue_r <= 16'b0001011110111011; rvalue_r <= 16'b0001011111001000;end
            11'b00111011111: begin lvalue_r <= 16'b0001011111001000; rvalue_r <= 16'b0001011111010101;end
            11'b00111100000: begin lvalue_r <= 16'b0001011111010101; rvalue_r <= 16'b0001011111100010;end
            11'b00111100001: begin lvalue_r <= 16'b0001011111100010; rvalue_r <= 16'b0001011111101111;end
            11'b00111100010: begin lvalue_r <= 16'b0001011111101111; rvalue_r <= 16'b0001011111111100;end
            11'b00111100011: begin lvalue_r <= 16'b0001011111111100; rvalue_r <= 16'b0001100000001001;end
            11'b00111100100: begin lvalue_r <= 16'b0001100000001001; rvalue_r <= 16'b0001100000010110;end
            11'b00111100101: begin lvalue_r <= 16'b0001100000010110; rvalue_r <= 16'b0001100000100011;end
            11'b00111100110: begin lvalue_r <= 16'b0001100000100011; rvalue_r <= 16'b0001100000110000;end
            11'b00111100111: begin lvalue_r <= 16'b0001100000110000; rvalue_r <= 16'b0001100000111101;end
            11'b00111101000: begin lvalue_r <= 16'b0001100000111101; rvalue_r <= 16'b0001100001001010;end
            11'b00111101001: begin lvalue_r <= 16'b0001100001001010; rvalue_r <= 16'b0001100001010111;end
            11'b00111101010: begin lvalue_r <= 16'b0001100001010111; rvalue_r <= 16'b0001100001100100;end
            11'b00111101011: begin lvalue_r <= 16'b0001100001100100; rvalue_r <= 16'b0001100001110001;end
            11'b00111101100: begin lvalue_r <= 16'b0001100001110001; rvalue_r <= 16'b0001100001111110;end
            11'b00111101101: begin lvalue_r <= 16'b0001100001111110; rvalue_r <= 16'b0001100010001011;end
            11'b00111101110: begin lvalue_r <= 16'b0001100010001011; rvalue_r <= 16'b0001100010011000;end
            11'b00111101111: begin lvalue_r <= 16'b0001100010011000; rvalue_r <= 16'b0001100010100101;end
            11'b00111110000: begin lvalue_r <= 16'b0001100010100101; rvalue_r <= 16'b0001100010110010;end
            11'b00111110001: begin lvalue_r <= 16'b0001100010110010; rvalue_r <= 16'b0001100010111111;end
            11'b00111110010: begin lvalue_r <= 16'b0001100010111111; rvalue_r <= 16'b0001100011001100;end
            11'b00111110011: begin lvalue_r <= 16'b0001100011001100; rvalue_r <= 16'b0001100011011001;end
            11'b00111110100: begin lvalue_r <= 16'b0001100011011001; rvalue_r <= 16'b0001100011100110;end
            11'b00111110101: begin lvalue_r <= 16'b0001100011100110; rvalue_r <= 16'b0001100011110011;end
            11'b00111110110: begin lvalue_r <= 16'b0001100011110011; rvalue_r <= 16'b0001100100000000;end
            11'b00111110111: begin lvalue_r <= 16'b0001100100000000; rvalue_r <= 16'b0001100100001110;end
            11'b00111111000: begin lvalue_r <= 16'b0001100100001110; rvalue_r <= 16'b0001100100011011;end
            11'b00111111001: begin lvalue_r <= 16'b0001100100011011; rvalue_r <= 16'b0001100100101000;end
            11'b00111111010: begin lvalue_r <= 16'b0001100100101000; rvalue_r <= 16'b0001100100110101;end
            11'b00111111011: begin lvalue_r <= 16'b0001100100110101; rvalue_r <= 16'b0001100101000010;end
            11'b00111111100: begin lvalue_r <= 16'b0001100101000010; rvalue_r <= 16'b0001100101001111;end
            11'b00111111101: begin lvalue_r <= 16'b0001100101001111; rvalue_r <= 16'b0001100101011100;end
            11'b00111111110: begin lvalue_r <= 16'b0001100101011100; rvalue_r <= 16'b0001100101101001;end
            11'b00111111111: begin lvalue_r <= 16'b0001100101101001; rvalue_r <= 16'b0001100101110110;end
            11'b01000000000: begin lvalue_r <= 16'b0001100101110110; rvalue_r <= 16'b0001100110000011;end
            11'b01000000001: begin lvalue_r <= 16'b0001100110000011; rvalue_r <= 16'b0001100110010000;end
            11'b01000000010: begin lvalue_r <= 16'b0001100110010000; rvalue_r <= 16'b0001100110011101;end
            11'b01000000011: begin lvalue_r <= 16'b0001100110011101; rvalue_r <= 16'b0001100110101010;end
            11'b01000000100: begin lvalue_r <= 16'b0001100110101010; rvalue_r <= 16'b0001100110110111;end
            11'b01000000101: begin lvalue_r <= 16'b0001100110110111; rvalue_r <= 16'b0001100111000100;end
            11'b01000000110: begin lvalue_r <= 16'b0001100111000100; rvalue_r <= 16'b0001100111010001;end
            11'b01000000111: begin lvalue_r <= 16'b0001100111010001; rvalue_r <= 16'b0001100111011111;end
            11'b01000001000: begin lvalue_r <= 16'b0001100111011111; rvalue_r <= 16'b0001100111101100;end
            11'b01000001001: begin lvalue_r <= 16'b0001100111101100; rvalue_r <= 16'b0001100111111001;end
            11'b01000001010: begin lvalue_r <= 16'b0001100111111001; rvalue_r <= 16'b0001101000000110;end
            11'b01000001011: begin lvalue_r <= 16'b0001101000000110; rvalue_r <= 16'b0001101000010011;end
            11'b01000001100: begin lvalue_r <= 16'b0001101000010011; rvalue_r <= 16'b0001101000100000;end
            11'b01000001101: begin lvalue_r <= 16'b0001101000100000; rvalue_r <= 16'b0001101000101101;end
            11'b01000001110: begin lvalue_r <= 16'b0001101000101101; rvalue_r <= 16'b0001101000111010;end
            11'b01000001111: begin lvalue_r <= 16'b0001101000111010; rvalue_r <= 16'b0001101001000111;end
            11'b01000010000: begin lvalue_r <= 16'b0001101001000111; rvalue_r <= 16'b0001101001010100;end
            11'b01000010001: begin lvalue_r <= 16'b0001101001010100; rvalue_r <= 16'b0001101001100001;end
            11'b01000010010: begin lvalue_r <= 16'b0001101001100001; rvalue_r <= 16'b0001101001101111;end
            11'b01000010011: begin lvalue_r <= 16'b0001101001101111; rvalue_r <= 16'b0001101001111100;end
            11'b01000010100: begin lvalue_r <= 16'b0001101001111100; rvalue_r <= 16'b0001101010001001;end
            11'b01000010101: begin lvalue_r <= 16'b0001101010001001; rvalue_r <= 16'b0001101010010110;end
            11'b01000010110: begin lvalue_r <= 16'b0001101010010110; rvalue_r <= 16'b0001101010100011;end
            11'b01000010111: begin lvalue_r <= 16'b0001101010100011; rvalue_r <= 16'b0001101010110000;end
            11'b01000011000: begin lvalue_r <= 16'b0001101010110000; rvalue_r <= 16'b0001101010111101;end
            11'b01000011001: begin lvalue_r <= 16'b0001101010111101; rvalue_r <= 16'b0001101011001010;end
            11'b01000011010: begin lvalue_r <= 16'b0001101011001010; rvalue_r <= 16'b0001101011010111;end
            11'b01000011011: begin lvalue_r <= 16'b0001101011010111; rvalue_r <= 16'b0001101011100101;end
            11'b01000011100: begin lvalue_r <= 16'b0001101011100101; rvalue_r <= 16'b0001101011110010;end
            11'b01000011101: begin lvalue_r <= 16'b0001101011110010; rvalue_r <= 16'b0001101011111111;end
            11'b01000011110: begin lvalue_r <= 16'b0001101011111111; rvalue_r <= 16'b0001101100001100;end
            11'b01000011111: begin lvalue_r <= 16'b0001101100001100; rvalue_r <= 16'b0001101100011001;end
            11'b01000100000: begin lvalue_r <= 16'b0001101100011001; rvalue_r <= 16'b0001101100100110;end
            11'b01000100001: begin lvalue_r <= 16'b0001101100100110; rvalue_r <= 16'b0001101100110011;end
            11'b01000100010: begin lvalue_r <= 16'b0001101100110011; rvalue_r <= 16'b0001101101000000;end
            11'b01000100011: begin lvalue_r <= 16'b0001101101000000; rvalue_r <= 16'b0001101101001110;end
            11'b01000100100: begin lvalue_r <= 16'b0001101101001110; rvalue_r <= 16'b0001101101011011;end
            11'b01000100101: begin lvalue_r <= 16'b0001101101011011; rvalue_r <= 16'b0001101101101000;end
            11'b01000100110: begin lvalue_r <= 16'b0001101101101000; rvalue_r <= 16'b0001101101110101;end
            11'b01000100111: begin lvalue_r <= 16'b0001101101110101; rvalue_r <= 16'b0001101110000010;end
            11'b01000101000: begin lvalue_r <= 16'b0001101110000010; rvalue_r <= 16'b0001101110001111;end
            11'b01000101001: begin lvalue_r <= 16'b0001101110001111; rvalue_r <= 16'b0001101110011100;end
            11'b01000101010: begin lvalue_r <= 16'b0001101110011100; rvalue_r <= 16'b0001101110101010;end
            11'b01000101011: begin lvalue_r <= 16'b0001101110101010; rvalue_r <= 16'b0001101110110111;end
            11'b01000101100: begin lvalue_r <= 16'b0001101110110111; rvalue_r <= 16'b0001101111000100;end
            11'b01000101101: begin lvalue_r <= 16'b0001101111000100; rvalue_r <= 16'b0001101111010001;end
            11'b01000101110: begin lvalue_r <= 16'b0001101111010001; rvalue_r <= 16'b0001101111011110;end
            11'b01000101111: begin lvalue_r <= 16'b0001101111011110; rvalue_r <= 16'b0001101111101011;end
            11'b01000110000: begin lvalue_r <= 16'b0001101111101011; rvalue_r <= 16'b0001101111111001;end
            11'b01000110001: begin lvalue_r <= 16'b0001101111111001; rvalue_r <= 16'b0001110000000110;end
            11'b01000110010: begin lvalue_r <= 16'b0001110000000110; rvalue_r <= 16'b0001110000010011;end
            11'b01000110011: begin lvalue_r <= 16'b0001110000010011; rvalue_r <= 16'b0001110000100000;end
            11'b01000110100: begin lvalue_r <= 16'b0001110000100000; rvalue_r <= 16'b0001110000101101;end
            11'b01000110101: begin lvalue_r <= 16'b0001110000101101; rvalue_r <= 16'b0001110000111010;end
            11'b01000110110: begin lvalue_r <= 16'b0001110000111010; rvalue_r <= 16'b0001110001001000;end
            11'b01000110111: begin lvalue_r <= 16'b0001110001001000; rvalue_r <= 16'b0001110001010101;end
            11'b01000111000: begin lvalue_r <= 16'b0001110001010101; rvalue_r <= 16'b0001110001100010;end
            11'b01000111001: begin lvalue_r <= 16'b0001110001100010; rvalue_r <= 16'b0001110001101111;end
            11'b01000111010: begin lvalue_r <= 16'b0001110001101111; rvalue_r <= 16'b0001110001111100;end
            11'b01000111011: begin lvalue_r <= 16'b0001110001111100; rvalue_r <= 16'b0001110010001010;end
            11'b01000111100: begin lvalue_r <= 16'b0001110010001010; rvalue_r <= 16'b0001110010010111;end
            11'b01000111101: begin lvalue_r <= 16'b0001110010010111; rvalue_r <= 16'b0001110010100100;end
            11'b01000111110: begin lvalue_r <= 16'b0001110010100100; rvalue_r <= 16'b0001110010110001;end
            11'b01000111111: begin lvalue_r <= 16'b0001110010110001; rvalue_r <= 16'b0001110010111110;end
            11'b01001000000: begin lvalue_r <= 16'b0001110010111110; rvalue_r <= 16'b0001110011001100;end
            11'b01001000001: begin lvalue_r <= 16'b0001110011001100; rvalue_r <= 16'b0001110011011001;end
            11'b01001000010: begin lvalue_r <= 16'b0001110011011001; rvalue_r <= 16'b0001110011100110;end
            11'b01001000011: begin lvalue_r <= 16'b0001110011100110; rvalue_r <= 16'b0001110011110011;end
            11'b01001000100: begin lvalue_r <= 16'b0001110011110011; rvalue_r <= 16'b0001110100000000;end
            11'b01001000101: begin lvalue_r <= 16'b0001110100000000; rvalue_r <= 16'b0001110100001110;end
            11'b01001000110: begin lvalue_r <= 16'b0001110100001110; rvalue_r <= 16'b0001110100011011;end
            11'b01001000111: begin lvalue_r <= 16'b0001110100011011; rvalue_r <= 16'b0001110100101000;end
            11'b01001001000: begin lvalue_r <= 16'b0001110100101000; rvalue_r <= 16'b0001110100110101;end
            11'b01001001001: begin lvalue_r <= 16'b0001110100110101; rvalue_r <= 16'b0001110101000010;end
            11'b01001001010: begin lvalue_r <= 16'b0001110101000010; rvalue_r <= 16'b0001110101010000;end
            11'b01001001011: begin lvalue_r <= 16'b0001110101010000; rvalue_r <= 16'b0001110101011101;end
            11'b01001001100: begin lvalue_r <= 16'b0001110101011101; rvalue_r <= 16'b0001110101101010;end
            11'b01001001101: begin lvalue_r <= 16'b0001110101101010; rvalue_r <= 16'b0001110101110111;end
            11'b01001001110: begin lvalue_r <= 16'b0001110101110111; rvalue_r <= 16'b0001110110000101;end
            11'b01001001111: begin lvalue_r <= 16'b0001110110000101; rvalue_r <= 16'b0001110110010010;end
            11'b01001010000: begin lvalue_r <= 16'b0001110110010010; rvalue_r <= 16'b0001110110011111;end
            11'b01001010001: begin lvalue_r <= 16'b0001110110011111; rvalue_r <= 16'b0001110110101100;end
            11'b01001010010: begin lvalue_r <= 16'b0001110110101100; rvalue_r <= 16'b0001110110111010;end
            11'b01001010011: begin lvalue_r <= 16'b0001110110111010; rvalue_r <= 16'b0001110111000111;end
            11'b01001010100: begin lvalue_r <= 16'b0001110111000111; rvalue_r <= 16'b0001110111010100;end
            11'b01001010101: begin lvalue_r <= 16'b0001110111010100; rvalue_r <= 16'b0001110111100001;end
            11'b01001010110: begin lvalue_r <= 16'b0001110111100001; rvalue_r <= 16'b0001110111101111;end
            11'b01001010111: begin lvalue_r <= 16'b0001110111101111; rvalue_r <= 16'b0001110111111100;end
            11'b01001011000: begin lvalue_r <= 16'b0001110111111100; rvalue_r <= 16'b0001111000001001;end
            11'b01001011001: begin lvalue_r <= 16'b0001111000001001; rvalue_r <= 16'b0001111000010110;end
            11'b01001011010: begin lvalue_r <= 16'b0001111000010110; rvalue_r <= 16'b0001111000100100;end
            11'b01001011011: begin lvalue_r <= 16'b0001111000100100; rvalue_r <= 16'b0001111000110001;end
            11'b01001011100: begin lvalue_r <= 16'b0001111000110001; rvalue_r <= 16'b0001111000111110;end
            11'b01001011101: begin lvalue_r <= 16'b0001111000111110; rvalue_r <= 16'b0001111001001011;end
            11'b01001011110: begin lvalue_r <= 16'b0001111001001011; rvalue_r <= 16'b0001111001011001;end
            11'b01001011111: begin lvalue_r <= 16'b0001111001011001; rvalue_r <= 16'b0001111001100110;end
            11'b01001100000: begin lvalue_r <= 16'b0001111001100110; rvalue_r <= 16'b0001111001110011;end
            11'b01001100001: begin lvalue_r <= 16'b0001111001110011; rvalue_r <= 16'b0001111010000000;end
            11'b01001100010: begin lvalue_r <= 16'b0001111010000000; rvalue_r <= 16'b0001111010001110;end
            11'b01001100011: begin lvalue_r <= 16'b0001111010001110; rvalue_r <= 16'b0001111010011011;end
            11'b01001100100: begin lvalue_r <= 16'b0001111010011011; rvalue_r <= 16'b0001111010101000;end
            11'b01001100101: begin lvalue_r <= 16'b0001111010101000; rvalue_r <= 16'b0001111010110110;end
            11'b01001100110: begin lvalue_r <= 16'b0001111010110110; rvalue_r <= 16'b0001111011000011;end
            11'b01001100111: begin lvalue_r <= 16'b0001111011000011; rvalue_r <= 16'b0001111011010000;end
            11'b01001101000: begin lvalue_r <= 16'b0001111011010000; rvalue_r <= 16'b0001111011011101;end
            11'b01001101001: begin lvalue_r <= 16'b0001111011011101; rvalue_r <= 16'b0001111011101011;end
            11'b01001101010: begin lvalue_r <= 16'b0001111011101011; rvalue_r <= 16'b0001111011111000;end
            11'b01001101011: begin lvalue_r <= 16'b0001111011111000; rvalue_r <= 16'b0001111100000101;end
            11'b01001101100: begin lvalue_r <= 16'b0001111100000101; rvalue_r <= 16'b0001111100010011;end
            11'b01001101101: begin lvalue_r <= 16'b0001111100010011; rvalue_r <= 16'b0001111100100000;end
            11'b01001101110: begin lvalue_r <= 16'b0001111100100000; rvalue_r <= 16'b0001111100101101;end
            11'b01001101111: begin lvalue_r <= 16'b0001111100101101; rvalue_r <= 16'b0001111100111011;end
            11'b01001110000: begin lvalue_r <= 16'b0001111100111011; rvalue_r <= 16'b0001111101001000;end
            11'b01001110001: begin lvalue_r <= 16'b0001111101001000; rvalue_r <= 16'b0001111101010101;end
            11'b01001110010: begin lvalue_r <= 16'b0001111101010101; rvalue_r <= 16'b0001111101100011;end
            11'b01001110011: begin lvalue_r <= 16'b0001111101100011; rvalue_r <= 16'b0001111101110000;end
            11'b01001110100: begin lvalue_r <= 16'b0001111101110000; rvalue_r <= 16'b0001111101111101;end
            11'b01001110101: begin lvalue_r <= 16'b0001111101111101; rvalue_r <= 16'b0001111110001011;end
            11'b01001110110: begin lvalue_r <= 16'b0001111110001011; rvalue_r <= 16'b0001111110011000;end
            11'b01001110111: begin lvalue_r <= 16'b0001111110011000; rvalue_r <= 16'b0001111110100101;end
            11'b01001111000: begin lvalue_r <= 16'b0001111110100101; rvalue_r <= 16'b0001111110110011;end
            11'b01001111001: begin lvalue_r <= 16'b0001111110110011; rvalue_r <= 16'b0001111111000000;end
            11'b01001111010: begin lvalue_r <= 16'b0001111111000000; rvalue_r <= 16'b0001111111001101;end
            11'b01001111011: begin lvalue_r <= 16'b0001111111001101; rvalue_r <= 16'b0001111111011011;end
            11'b01001111100: begin lvalue_r <= 16'b0001111111011011; rvalue_r <= 16'b0001111111101000;end
            11'b01001111101: begin lvalue_r <= 16'b0001111111101000; rvalue_r <= 16'b0001111111110101;end
            11'b01001111110: begin lvalue_r <= 16'b0001111111110101; rvalue_r <= 16'b0010000000000011;end
            11'b01001111111: begin lvalue_r <= 16'b0010000000000011; rvalue_r <= 16'b0010000000010000;end
            11'b01010000000: begin lvalue_r <= 16'b0010000000010000; rvalue_r <= 16'b0010000000011101;end
            11'b01010000001: begin lvalue_r <= 16'b0010000000011101; rvalue_r <= 16'b0010000000101011;end
            11'b01010000010: begin lvalue_r <= 16'b0010000000101011; rvalue_r <= 16'b0010000000111000;end
            11'b01010000011: begin lvalue_r <= 16'b0010000000111000; rvalue_r <= 16'b0010000001000101;end
            11'b01010000100: begin lvalue_r <= 16'b0010000001000101; rvalue_r <= 16'b0010000001010011;end
            11'b01010000101: begin lvalue_r <= 16'b0010000001010011; rvalue_r <= 16'b0010000001100000;end
            11'b01010000110: begin lvalue_r <= 16'b0010000001100000; rvalue_r <= 16'b0010000001101110;end
            11'b01010000111: begin lvalue_r <= 16'b0010000001101110; rvalue_r <= 16'b0010000001111011;end
            11'b01010001000: begin lvalue_r <= 16'b0010000001111011; rvalue_r <= 16'b0010000010001000;end
            11'b01010001001: begin lvalue_r <= 16'b0010000010001000; rvalue_r <= 16'b0010000010010110;end
            11'b01010001010: begin lvalue_r <= 16'b0010000010010110; rvalue_r <= 16'b0010000010100011;end
            11'b01010001011: begin lvalue_r <= 16'b0010000010100011; rvalue_r <= 16'b0010000010110000;end
            11'b01010001100: begin lvalue_r <= 16'b0010000010110000; rvalue_r <= 16'b0010000010111110;end
            11'b01010001101: begin lvalue_r <= 16'b0010000010111110; rvalue_r <= 16'b0010000011001011;end
            11'b01010001110: begin lvalue_r <= 16'b0010000011001011; rvalue_r <= 16'b0010000011011001;end
            11'b01010001111: begin lvalue_r <= 16'b0010000011011001; rvalue_r <= 16'b0010000011100110;end
            11'b01010010000: begin lvalue_r <= 16'b0010000011100110; rvalue_r <= 16'b0010000011110011;end
            11'b01010010001: begin lvalue_r <= 16'b0010000011110011; rvalue_r <= 16'b0010000100000001;end
            11'b01010010010: begin lvalue_r <= 16'b0010000100000001; rvalue_r <= 16'b0010000100001110;end
            11'b01010010011: begin lvalue_r <= 16'b0010000100001110; rvalue_r <= 16'b0010000100011100;end
            11'b01010010100: begin lvalue_r <= 16'b0010000100011100; rvalue_r <= 16'b0010000100101001;end
            11'b01010010101: begin lvalue_r <= 16'b0010000100101001; rvalue_r <= 16'b0010000100110110;end
            11'b01010010110: begin lvalue_r <= 16'b0010000100110110; rvalue_r <= 16'b0010000101000100;end
            11'b01010010111: begin lvalue_r <= 16'b0010000101000100; rvalue_r <= 16'b0010000101010001;end
            11'b01010011000: begin lvalue_r <= 16'b0010000101010001; rvalue_r <= 16'b0010000101011111;end
            11'b01010011001: begin lvalue_r <= 16'b0010000101011111; rvalue_r <= 16'b0010000101101100;end
            11'b01010011010: begin lvalue_r <= 16'b0010000101101100; rvalue_r <= 16'b0010000101111001;end
            11'b01010011011: begin lvalue_r <= 16'b0010000101111001; rvalue_r <= 16'b0010000110000111;end
            11'b01010011100: begin lvalue_r <= 16'b0010000110000111; rvalue_r <= 16'b0010000110010100;end
            11'b01010011101: begin lvalue_r <= 16'b0010000110010100; rvalue_r <= 16'b0010000110100010;end
            11'b01010011110: begin lvalue_r <= 16'b0010000110100010; rvalue_r <= 16'b0010000110101111;end
            11'b01010011111: begin lvalue_r <= 16'b0010000110101111; rvalue_r <= 16'b0010000110111101;end
            11'b01010100000: begin lvalue_r <= 16'b0010000110111101; rvalue_r <= 16'b0010000111001010;end
            11'b01010100001: begin lvalue_r <= 16'b0010000111001010; rvalue_r <= 16'b0010000111011000;end
            11'b01010100010: begin lvalue_r <= 16'b0010000111011000; rvalue_r <= 16'b0010000111100101;end
            11'b01010100011: begin lvalue_r <= 16'b0010000111100101; rvalue_r <= 16'b0010000111110010;end
            11'b01010100100: begin lvalue_r <= 16'b0010000111110010; rvalue_r <= 16'b0010001000000000;end
            11'b01010100101: begin lvalue_r <= 16'b0010001000000000; rvalue_r <= 16'b0010001000001101;end
            11'b01010100110: begin lvalue_r <= 16'b0010001000001101; rvalue_r <= 16'b0010001000011011;end
            11'b01010100111: begin lvalue_r <= 16'b0010001000011011; rvalue_r <= 16'b0010001000101000;end
            11'b01010101000: begin lvalue_r <= 16'b0010001000101000; rvalue_r <= 16'b0010001000110110;end
            11'b01010101001: begin lvalue_r <= 16'b0010001000110110; rvalue_r <= 16'b0010001001000011;end
            11'b01010101010: begin lvalue_r <= 16'b0010001001000011; rvalue_r <= 16'b0010001001010001;end
            11'b01010101011: begin lvalue_r <= 16'b0010001001010001; rvalue_r <= 16'b0010001001011110;end
            11'b01010101100: begin lvalue_r <= 16'b0010001001011110; rvalue_r <= 16'b0010001001101100;end
            11'b01010101101: begin lvalue_r <= 16'b0010001001101100; rvalue_r <= 16'b0010001001111001;end
            11'b01010101110: begin lvalue_r <= 16'b0010001001111001; rvalue_r <= 16'b0010001010000111;end
            11'b01010101111: begin lvalue_r <= 16'b0010001010000111; rvalue_r <= 16'b0010001010010100;end
            11'b01010110000: begin lvalue_r <= 16'b0010001010010100; rvalue_r <= 16'b0010001010100010;end
            11'b01010110001: begin lvalue_r <= 16'b0010001010100010; rvalue_r <= 16'b0010001010101111;end
            11'b01010110010: begin lvalue_r <= 16'b0010001010101111; rvalue_r <= 16'b0010001010111100;end
            11'b01010110011: begin lvalue_r <= 16'b0010001010111100; rvalue_r <= 16'b0010001011001010;end
            11'b01010110100: begin lvalue_r <= 16'b0010001011001010; rvalue_r <= 16'b0010001011010111;end
            11'b01010110101: begin lvalue_r <= 16'b0010001011010111; rvalue_r <= 16'b0010001011100101;end
            11'b01010110110: begin lvalue_r <= 16'b0010001011100101; rvalue_r <= 16'b0010001011110010;end
            11'b01010110111: begin lvalue_r <= 16'b0010001011110010; rvalue_r <= 16'b0010001100000000;end
            11'b01010111000: begin lvalue_r <= 16'b0010001100000000; rvalue_r <= 16'b0010001100001101;end
            11'b01010111001: begin lvalue_r <= 16'b0010001100001101; rvalue_r <= 16'b0010001100011011;end
            11'b01010111010: begin lvalue_r <= 16'b0010001100011011; rvalue_r <= 16'b0010001100101001;end
            11'b01010111011: begin lvalue_r <= 16'b0010001100101001; rvalue_r <= 16'b0010001100110110;end
            11'b01010111100: begin lvalue_r <= 16'b0010001100110110; rvalue_r <= 16'b0010001101000100;end
            11'b01010111101: begin lvalue_r <= 16'b0010001101000100; rvalue_r <= 16'b0010001101010001;end
            11'b01010111110: begin lvalue_r <= 16'b0010001101010001; rvalue_r <= 16'b0010001101011111;end
            11'b01010111111: begin lvalue_r <= 16'b0010001101011111; rvalue_r <= 16'b0010001101101100;end
            11'b01011000000: begin lvalue_r <= 16'b0010001101101100; rvalue_r <= 16'b0010001101111010;end
            11'b01011000001: begin lvalue_r <= 16'b0010001101111010; rvalue_r <= 16'b0010001110000111;end
            11'b01011000010: begin lvalue_r <= 16'b0010001110000111; rvalue_r <= 16'b0010001110010101;end
            11'b01011000011: begin lvalue_r <= 16'b0010001110010101; rvalue_r <= 16'b0010001110100010;end
            11'b01011000100: begin lvalue_r <= 16'b0010001110100010; rvalue_r <= 16'b0010001110110000;end
            11'b01011000101: begin lvalue_r <= 16'b0010001110110000; rvalue_r <= 16'b0010001110111101;end
            11'b01011000110: begin lvalue_r <= 16'b0010001110111101; rvalue_r <= 16'b0010001111001011;end
            11'b01011000111: begin lvalue_r <= 16'b0010001111001011; rvalue_r <= 16'b0010001111011000;end
            11'b01011001000: begin lvalue_r <= 16'b0010001111011000; rvalue_r <= 16'b0010001111100110;end
            11'b01011001001: begin lvalue_r <= 16'b0010001111100110; rvalue_r <= 16'b0010001111110100;end
            11'b01011001010: begin lvalue_r <= 16'b0010001111110100; rvalue_r <= 16'b0010010000000001;end
            11'b01011001011: begin lvalue_r <= 16'b0010010000000001; rvalue_r <= 16'b0010010000001111;end
            11'b01011001100: begin lvalue_r <= 16'b0010010000001111; rvalue_r <= 16'b0010010000011100;end
            11'b01011001101: begin lvalue_r <= 16'b0010010000011100; rvalue_r <= 16'b0010010000101010;end
            11'b01011001110: begin lvalue_r <= 16'b0010010000101010; rvalue_r <= 16'b0010010000110111;end
            11'b01011001111: begin lvalue_r <= 16'b0010010000110111; rvalue_r <= 16'b0010010001000101;end
            11'b01011010000: begin lvalue_r <= 16'b0010010001000101; rvalue_r <= 16'b0010010001010011;end
            11'b01011010001: begin lvalue_r <= 16'b0010010001010011; rvalue_r <= 16'b0010010001100000;end
            11'b01011010010: begin lvalue_r <= 16'b0010010001100000; rvalue_r <= 16'b0010010001101110;end
            11'b01011010011: begin lvalue_r <= 16'b0010010001101110; rvalue_r <= 16'b0010010001111011;end
            11'b01011010100: begin lvalue_r <= 16'b0010010001111011; rvalue_r <= 16'b0010010010001001;end
            11'b01011010101: begin lvalue_r <= 16'b0010010010001001; rvalue_r <= 16'b0010010010010110;end
            11'b01011010110: begin lvalue_r <= 16'b0010010010010110; rvalue_r <= 16'b0010010010100100;end
            11'b01011010111: begin lvalue_r <= 16'b0010010010100100; rvalue_r <= 16'b0010010010110010;end
            11'b01011011000: begin lvalue_r <= 16'b0010010010110010; rvalue_r <= 16'b0010010010111111;end
            11'b01011011001: begin lvalue_r <= 16'b0010010010111111; rvalue_r <= 16'b0010010011001101;end
            11'b01011011010: begin lvalue_r <= 16'b0010010011001101; rvalue_r <= 16'b0010010011011010;end
            11'b01011011011: begin lvalue_r <= 16'b0010010011011010; rvalue_r <= 16'b0010010011101000;end
            11'b01011011100: begin lvalue_r <= 16'b0010010011101000; rvalue_r <= 16'b0010010011110110;end
            11'b01011011101: begin lvalue_r <= 16'b0010010011110110; rvalue_r <= 16'b0010010100000011;end
            11'b01011011110: begin lvalue_r <= 16'b0010010100000011; rvalue_r <= 16'b0010010100010001;end
            11'b01011011111: begin lvalue_r <= 16'b0010010100010001; rvalue_r <= 16'b0010010100011111;end
            11'b01011100000: begin lvalue_r <= 16'b0010010100011111; rvalue_r <= 16'b0010010100101100;end
            11'b01011100001: begin lvalue_r <= 16'b0010010100101100; rvalue_r <= 16'b0010010100111010;end
            11'b01011100010: begin lvalue_r <= 16'b0010010100111010; rvalue_r <= 16'b0010010101000111;end
            11'b01011100011: begin lvalue_r <= 16'b0010010101000111; rvalue_r <= 16'b0010010101010101;end
            11'b01011100100: begin lvalue_r <= 16'b0010010101010101; rvalue_r <= 16'b0010010101100011;end
            11'b01011100101: begin lvalue_r <= 16'b0010010101100011; rvalue_r <= 16'b0010010101110000;end
            11'b01011100110: begin lvalue_r <= 16'b0010010101110000; rvalue_r <= 16'b0010010101111110;end
            11'b01011100111: begin lvalue_r <= 16'b0010010101111110; rvalue_r <= 16'b0010010110001100;end
            11'b01011101000: begin lvalue_r <= 16'b0010010110001100; rvalue_r <= 16'b0010010110011001;end
            11'b01011101001: begin lvalue_r <= 16'b0010010110011001; rvalue_r <= 16'b0010010110100111;end
            11'b01011101010: begin lvalue_r <= 16'b0010010110100111; rvalue_r <= 16'b0010010110110101;end
            11'b01011101011: begin lvalue_r <= 16'b0010010110110101; rvalue_r <= 16'b0010010111000010;end
            11'b01011101100: begin lvalue_r <= 16'b0010010111000010; rvalue_r <= 16'b0010010111010000;end
            11'b01011101101: begin lvalue_r <= 16'b0010010111010000; rvalue_r <= 16'b0010010111011110;end
            11'b01011101110: begin lvalue_r <= 16'b0010010111011110; rvalue_r <= 16'b0010010111101011;end
            11'b01011101111: begin lvalue_r <= 16'b0010010111101011; rvalue_r <= 16'b0010010111111001;end
            11'b01011110000: begin lvalue_r <= 16'b0010010111111001; rvalue_r <= 16'b0010011000000111;end
            11'b01011110001: begin lvalue_r <= 16'b0010011000000111; rvalue_r <= 16'b0010011000010100;end
            11'b01011110010: begin lvalue_r <= 16'b0010011000010100; rvalue_r <= 16'b0010011000100010;end
            11'b01011110011: begin lvalue_r <= 16'b0010011000100010; rvalue_r <= 16'b0010011000110000;end
            11'b01011110100: begin lvalue_r <= 16'b0010011000110000; rvalue_r <= 16'b0010011000111101;end
            11'b01011110101: begin lvalue_r <= 16'b0010011000111101; rvalue_r <= 16'b0010011001001011;end
            11'b01011110110: begin lvalue_r <= 16'b0010011001001011; rvalue_r <= 16'b0010011001011001;end
            11'b01011110111: begin lvalue_r <= 16'b0010011001011001; rvalue_r <= 16'b0010011001100110;end
            11'b01011111000: begin lvalue_r <= 16'b0010011001100110; rvalue_r <= 16'b0010011001110100;end
            11'b01011111001: begin lvalue_r <= 16'b0010011001110100; rvalue_r <= 16'b0010011010000010;end
            11'b01011111010: begin lvalue_r <= 16'b0010011010000010; rvalue_r <= 16'b0010011010001111;end
            11'b01011111011: begin lvalue_r <= 16'b0010011010001111; rvalue_r <= 16'b0010011010011101;end
            11'b01011111100: begin lvalue_r <= 16'b0010011010011101; rvalue_r <= 16'b0010011010101011;end
            11'b01011111101: begin lvalue_r <= 16'b0010011010101011; rvalue_r <= 16'b0010011010111001;end
            11'b01011111110: begin lvalue_r <= 16'b0010011010111001; rvalue_r <= 16'b0010011011000110;end
            11'b01011111111: begin lvalue_r <= 16'b0010011011000110; rvalue_r <= 16'b0010011011010100;end
            11'b01100000000: begin lvalue_r <= 16'b0010011011010100; rvalue_r <= 16'b0010011011100010;end
            11'b01100000001: begin lvalue_r <= 16'b0010011011100010; rvalue_r <= 16'b0010011011110000;end
            11'b01100000010: begin lvalue_r <= 16'b0010011011110000; rvalue_r <= 16'b0010011011111101;end
            11'b01100000011: begin lvalue_r <= 16'b0010011011111101; rvalue_r <= 16'b0010011100001011;end
            11'b01100000100: begin lvalue_r <= 16'b0010011100001011; rvalue_r <= 16'b0010011100011001;end
            11'b01100000101: begin lvalue_r <= 16'b0010011100011001; rvalue_r <= 16'b0010011100100110;end
            11'b01100000110: begin lvalue_r <= 16'b0010011100100110; rvalue_r <= 16'b0010011100110100;end
            11'b01100000111: begin lvalue_r <= 16'b0010011100110100; rvalue_r <= 16'b0010011101000010;end
            11'b01100001000: begin lvalue_r <= 16'b0010011101000010; rvalue_r <= 16'b0010011101010000;end
            11'b01100001001: begin lvalue_r <= 16'b0010011101010000; rvalue_r <= 16'b0010011101011101;end
            11'b01100001010: begin lvalue_r <= 16'b0010011101011101; rvalue_r <= 16'b0010011101101011;end
            11'b01100001011: begin lvalue_r <= 16'b0010011101101011; rvalue_r <= 16'b0010011101111001;end
            11'b01100001100: begin lvalue_r <= 16'b0010011101111001; rvalue_r <= 16'b0010011110000111;end
            11'b01100001101: begin lvalue_r <= 16'b0010011110000111; rvalue_r <= 16'b0010011110010100;end
            11'b01100001110: begin lvalue_r <= 16'b0010011110010100; rvalue_r <= 16'b0010011110100010;end
            11'b01100001111: begin lvalue_r <= 16'b0010011110100010; rvalue_r <= 16'b0010011110110000;end
            11'b01100010000: begin lvalue_r <= 16'b0010011110110000; rvalue_r <= 16'b0010011110111110;end
            11'b01100010001: begin lvalue_r <= 16'b0010011110111110; rvalue_r <= 16'b0010011111001100;end
            11'b01100010010: begin lvalue_r <= 16'b0010011111001100; rvalue_r <= 16'b0010011111011001;end
            11'b01100010011: begin lvalue_r <= 16'b0010011111011001; rvalue_r <= 16'b0010011111100111;end
            11'b01100010100: begin lvalue_r <= 16'b0010011111100111; rvalue_r <= 16'b0010011111110101;end
            11'b01100010101: begin lvalue_r <= 16'b0010011111110101; rvalue_r <= 16'b0010100000000011;end
            11'b01100010110: begin lvalue_r <= 16'b0010100000000011; rvalue_r <= 16'b0010100000010001;end
            11'b01100010111: begin lvalue_r <= 16'b0010100000010001; rvalue_r <= 16'b0010100000011110;end
            11'b01100011000: begin lvalue_r <= 16'b0010100000011110; rvalue_r <= 16'b0010100000101100;end
            11'b01100011001: begin lvalue_r <= 16'b0010100000101100; rvalue_r <= 16'b0010100000111010;end
            11'b01100011010: begin lvalue_r <= 16'b0010100000111010; rvalue_r <= 16'b0010100001001000;end
            11'b01100011011: begin lvalue_r <= 16'b0010100001001000; rvalue_r <= 16'b0010100001010110;end
            11'b01100011100: begin lvalue_r <= 16'b0010100001010110; rvalue_r <= 16'b0010100001100011;end
            11'b01100011101: begin lvalue_r <= 16'b0010100001100011; rvalue_r <= 16'b0010100001110001;end
            11'b01100011110: begin lvalue_r <= 16'b0010100001110001; rvalue_r <= 16'b0010100001111111;end
            11'b01100011111: begin lvalue_r <= 16'b0010100001111111; rvalue_r <= 16'b0010100010001101;end
            11'b01100100000: begin lvalue_r <= 16'b0010100010001101; rvalue_r <= 16'b0010100010011011;end
            11'b01100100001: begin lvalue_r <= 16'b0010100010011011; rvalue_r <= 16'b0010100010101001;end
            11'b01100100010: begin lvalue_r <= 16'b0010100010101001; rvalue_r <= 16'b0010100010110110;end
            11'b01100100011: begin lvalue_r <= 16'b0010100010110110; rvalue_r <= 16'b0010100011000100;end
            11'b01100100100: begin lvalue_r <= 16'b0010100011000100; rvalue_r <= 16'b0010100011010010;end
            11'b01100100101: begin lvalue_r <= 16'b0010100011010010; rvalue_r <= 16'b0010100011100000;end
            11'b01100100110: begin lvalue_r <= 16'b0010100011100000; rvalue_r <= 16'b0010100011101110;end
            11'b01100100111: begin lvalue_r <= 16'b0010100011101110; rvalue_r <= 16'b0010100011111100;end
            11'b01100101000: begin lvalue_r <= 16'b0010100011111100; rvalue_r <= 16'b0010100100001001;end
            11'b01100101001: begin lvalue_r <= 16'b0010100100001001; rvalue_r <= 16'b0010100100010111;end
            11'b01100101010: begin lvalue_r <= 16'b0010100100010111; rvalue_r <= 16'b0010100100100101;end
            11'b01100101011: begin lvalue_r <= 16'b0010100100100101; rvalue_r <= 16'b0010100100110011;end
            11'b01100101100: begin lvalue_r <= 16'b0010100100110011; rvalue_r <= 16'b0010100101000001;end
            11'b01100101101: begin lvalue_r <= 16'b0010100101000001; rvalue_r <= 16'b0010100101001111;end
            11'b01100101110: begin lvalue_r <= 16'b0010100101001111; rvalue_r <= 16'b0010100101011101;end
            11'b01100101111: begin lvalue_r <= 16'b0010100101011101; rvalue_r <= 16'b0010100101101011;end
            11'b01100110000: begin lvalue_r <= 16'b0010100101101011; rvalue_r <= 16'b0010100101111000;end
            11'b01100110001: begin lvalue_r <= 16'b0010100101111000; rvalue_r <= 16'b0010100110000110;end
            11'b01100110010: begin lvalue_r <= 16'b0010100110000110; rvalue_r <= 16'b0010100110010100;end
            11'b01100110011: begin lvalue_r <= 16'b0010100110010100; rvalue_r <= 16'b0010100110100010;end
            11'b01100110100: begin lvalue_r <= 16'b0010100110100010; rvalue_r <= 16'b0010100110110000;end
            11'b01100110101: begin lvalue_r <= 16'b0010100110110000; rvalue_r <= 16'b0010100110111110;end
            11'b01100110110: begin lvalue_r <= 16'b0010100110111110; rvalue_r <= 16'b0010100111001100;end
            11'b01100110111: begin lvalue_r <= 16'b0010100111001100; rvalue_r <= 16'b0010100111011010;end
            11'b01100111000: begin lvalue_r <= 16'b0010100111011010; rvalue_r <= 16'b0010100111101000;end
            11'b01100111001: begin lvalue_r <= 16'b0010100111101000; rvalue_r <= 16'b0010100111110110;end
            11'b01100111010: begin lvalue_r <= 16'b0010100111110110; rvalue_r <= 16'b0010101000000011;end
            11'b01100111011: begin lvalue_r <= 16'b0010101000000011; rvalue_r <= 16'b0010101000010001;end
            11'b01100111100: begin lvalue_r <= 16'b0010101000010001; rvalue_r <= 16'b0010101000011111;end
            11'b01100111101: begin lvalue_r <= 16'b0010101000011111; rvalue_r <= 16'b0010101000101101;end
            11'b01100111110: begin lvalue_r <= 16'b0010101000101101; rvalue_r <= 16'b0010101000111011;end
            11'b01100111111: begin lvalue_r <= 16'b0010101000111011; rvalue_r <= 16'b0010101001001001;end
            11'b01101000000: begin lvalue_r <= 16'b0010101001001001; rvalue_r <= 16'b0010101001010111;end
            11'b01101000001: begin lvalue_r <= 16'b0010101001010111; rvalue_r <= 16'b0010101001100101;end
            11'b01101000010: begin lvalue_r <= 16'b0010101001100101; rvalue_r <= 16'b0010101001110011;end
            11'b01101000011: begin lvalue_r <= 16'b0010101001110011; rvalue_r <= 16'b0010101010000001;end
            11'b01101000100: begin lvalue_r <= 16'b0010101010000001; rvalue_r <= 16'b0010101010001111;end
            11'b01101000101: begin lvalue_r <= 16'b0010101010001111; rvalue_r <= 16'b0010101010011101;end
            11'b01101000110: begin lvalue_r <= 16'b0010101010011101; rvalue_r <= 16'b0010101010101011;end
            11'b01101000111: begin lvalue_r <= 16'b0010101010101011; rvalue_r <= 16'b0010101010111001;end
            11'b01101001000: begin lvalue_r <= 16'b0010101010111001; rvalue_r <= 16'b0010101011000111;end
            11'b01101001001: begin lvalue_r <= 16'b0010101011000111; rvalue_r <= 16'b0010101011010101;end
            11'b01101001010: begin lvalue_r <= 16'b0010101011010101; rvalue_r <= 16'b0010101011100011;end
            11'b01101001011: begin lvalue_r <= 16'b0010101011100011; rvalue_r <= 16'b0010101011110001;end
            11'b01101001100: begin lvalue_r <= 16'b0010101011110001; rvalue_r <= 16'b0010101011111111;end
            11'b01101001101: begin lvalue_r <= 16'b0010101011111111; rvalue_r <= 16'b0010101100001101;end
            11'b01101001110: begin lvalue_r <= 16'b0010101100001101; rvalue_r <= 16'b0010101100011011;end
            11'b01101001111: begin lvalue_r <= 16'b0010101100011011; rvalue_r <= 16'b0010101100101001;end
            11'b01101010000: begin lvalue_r <= 16'b0010101100101001; rvalue_r <= 16'b0010101100110111;end
            11'b01101010001: begin lvalue_r <= 16'b0010101100110111; rvalue_r <= 16'b0010101101000101;end
            11'b01101010010: begin lvalue_r <= 16'b0010101101000101; rvalue_r <= 16'b0010101101010011;end
            11'b01101010011: begin lvalue_r <= 16'b0010101101010011; rvalue_r <= 16'b0010101101100001;end
            11'b01101010100: begin lvalue_r <= 16'b0010101101100001; rvalue_r <= 16'b0010101101101111;end
            11'b01101010101: begin lvalue_r <= 16'b0010101101101111; rvalue_r <= 16'b0010101101111101;end
            11'b01101010110: begin lvalue_r <= 16'b0010101101111101; rvalue_r <= 16'b0010101110001011;end
            11'b01101010111: begin lvalue_r <= 16'b0010101110001011; rvalue_r <= 16'b0010101110011001;end
            11'b01101011000: begin lvalue_r <= 16'b0010101110011001; rvalue_r <= 16'b0010101110100111;end
            11'b01101011001: begin lvalue_r <= 16'b0010101110100111; rvalue_r <= 16'b0010101110110101;end
            11'b01101011010: begin lvalue_r <= 16'b0010101110110101; rvalue_r <= 16'b0010101111000011;end
            11'b01101011011: begin lvalue_r <= 16'b0010101111000011; rvalue_r <= 16'b0010101111010001;end
            11'b01101011100: begin lvalue_r <= 16'b0010101111010001; rvalue_r <= 16'b0010101111011111;end
            11'b01101011101: begin lvalue_r <= 16'b0010101111011111; rvalue_r <= 16'b0010101111101101;end
            11'b01101011110: begin lvalue_r <= 16'b0010101111101101; rvalue_r <= 16'b0010101111111011;end
            11'b01101011111: begin lvalue_r <= 16'b0010101111111011; rvalue_r <= 16'b0010110000001001;end
            11'b01101100000: begin lvalue_r <= 16'b0010110000001001; rvalue_r <= 16'b0010110000010111;end
            11'b01101100001: begin lvalue_r <= 16'b0010110000010111; rvalue_r <= 16'b0010110000100101;end
            11'b01101100010: begin lvalue_r <= 16'b0010110000100101; rvalue_r <= 16'b0010110000110011;end
            11'b01101100011: begin lvalue_r <= 16'b0010110000110011; rvalue_r <= 16'b0010110001000001;end
            11'b01101100100: begin lvalue_r <= 16'b0010110001000001; rvalue_r <= 16'b0010110001001111;end
            11'b01101100101: begin lvalue_r <= 16'b0010110001001111; rvalue_r <= 16'b0010110001011101;end
            11'b01101100110: begin lvalue_r <= 16'b0010110001011101; rvalue_r <= 16'b0010110001101011;end
            11'b01101100111: begin lvalue_r <= 16'b0010110001101011; rvalue_r <= 16'b0010110001111001;end
            11'b01101101000: begin lvalue_r <= 16'b0010110001111001; rvalue_r <= 16'b0010110010001000;end
            11'b01101101001: begin lvalue_r <= 16'b0010110010001000; rvalue_r <= 16'b0010110010010110;end
            11'b01101101010: begin lvalue_r <= 16'b0010110010010110; rvalue_r <= 16'b0010110010100100;end
            11'b01101101011: begin lvalue_r <= 16'b0010110010100100; rvalue_r <= 16'b0010110010110010;end
            11'b01101101100: begin lvalue_r <= 16'b0010110010110010; rvalue_r <= 16'b0010110011000000;end
            11'b01101101101: begin lvalue_r <= 16'b0010110011000000; rvalue_r <= 16'b0010110011001110;end
            11'b01101101110: begin lvalue_r <= 16'b0010110011001110; rvalue_r <= 16'b0010110011011100;end
            11'b01101101111: begin lvalue_r <= 16'b0010110011011100; rvalue_r <= 16'b0010110011101010;end
            11'b01101110000: begin lvalue_r <= 16'b0010110011101010; rvalue_r <= 16'b0010110011111000;end
            11'b01101110001: begin lvalue_r <= 16'b0010110011111000; rvalue_r <= 16'b0010110100000111;end
            11'b01101110010: begin lvalue_r <= 16'b0010110100000111; rvalue_r <= 16'b0010110100010101;end
            11'b01101110011: begin lvalue_r <= 16'b0010110100010101; rvalue_r <= 16'b0010110100100011;end
            11'b01101110100: begin lvalue_r <= 16'b0010110100100011; rvalue_r <= 16'b0010110100110001;end
            11'b01101110101: begin lvalue_r <= 16'b0010110100110001; rvalue_r <= 16'b0010110100111111;end
            11'b01101110110: begin lvalue_r <= 16'b0010110100111111; rvalue_r <= 16'b0010110101001101;end
            11'b01101110111: begin lvalue_r <= 16'b0010110101001101; rvalue_r <= 16'b0010110101011011;end
            11'b01101111000: begin lvalue_r <= 16'b0010110101011011; rvalue_r <= 16'b0010110101101001;end
            11'b01101111001: begin lvalue_r <= 16'b0010110101101001; rvalue_r <= 16'b0010110101111000;end
            11'b01101111010: begin lvalue_r <= 16'b0010110101111000; rvalue_r <= 16'b0010110110000110;end
            11'b01101111011: begin lvalue_r <= 16'b0010110110000110; rvalue_r <= 16'b0010110110010100;end
            11'b01101111100: begin lvalue_r <= 16'b0010110110010100; rvalue_r <= 16'b0010110110100010;end
            11'b01101111101: begin lvalue_r <= 16'b0010110110100010; rvalue_r <= 16'b0010110110110000;end
            11'b01101111110: begin lvalue_r <= 16'b0010110110110000; rvalue_r <= 16'b0010110110111110;end
            11'b01101111111: begin lvalue_r <= 16'b0010110110111110; rvalue_r <= 16'b0010110111001101;end
            11'b01110000000: begin lvalue_r <= 16'b0010110111001101; rvalue_r <= 16'b0010110111011011;end
            11'b01110000001: begin lvalue_r <= 16'b0010110111011011; rvalue_r <= 16'b0010110111101001;end
            11'b01110000010: begin lvalue_r <= 16'b0010110111101001; rvalue_r <= 16'b0010110111110111;end
            11'b01110000011: begin lvalue_r <= 16'b0010110111110111; rvalue_r <= 16'b0010111000000101;end
            11'b01110000100: begin lvalue_r <= 16'b0010111000000101; rvalue_r <= 16'b0010111000010100;end
            11'b01110000101: begin lvalue_r <= 16'b0010111000010100; rvalue_r <= 16'b0010111000100010;end
            11'b01110000110: begin lvalue_r <= 16'b0010111000100010; rvalue_r <= 16'b0010111000110000;end
            11'b01110000111: begin lvalue_r <= 16'b0010111000110000; rvalue_r <= 16'b0010111000111110;end
            11'b01110001000: begin lvalue_r <= 16'b0010111000111110; rvalue_r <= 16'b0010111001001100;end
            11'b01110001001: begin lvalue_r <= 16'b0010111001001100; rvalue_r <= 16'b0010111001011011;end
            11'b01110001010: begin lvalue_r <= 16'b0010111001011011; rvalue_r <= 16'b0010111001101001;end
            11'b01110001011: begin lvalue_r <= 16'b0010111001101001; rvalue_r <= 16'b0010111001110111;end
            11'b01110001100: begin lvalue_r <= 16'b0010111001110111; rvalue_r <= 16'b0010111010000101;end
            11'b01110001101: begin lvalue_r <= 16'b0010111010000101; rvalue_r <= 16'b0010111010010011;end
            11'b01110001110: begin lvalue_r <= 16'b0010111010010011; rvalue_r <= 16'b0010111010100010;end
            11'b01110001111: begin lvalue_r <= 16'b0010111010100010; rvalue_r <= 16'b0010111010110000;end
            11'b01110010000: begin lvalue_r <= 16'b0010111010110000; rvalue_r <= 16'b0010111010111110;end
            11'b01110010001: begin lvalue_r <= 16'b0010111010111110; rvalue_r <= 16'b0010111011001100;end
            11'b01110010010: begin lvalue_r <= 16'b0010111011001100; rvalue_r <= 16'b0010111011011011;end
            11'b01110010011: begin lvalue_r <= 16'b0010111011011011; rvalue_r <= 16'b0010111011101001;end
            11'b01110010100: begin lvalue_r <= 16'b0010111011101001; rvalue_r <= 16'b0010111011110111;end
            11'b01110010101: begin lvalue_r <= 16'b0010111011110111; rvalue_r <= 16'b0010111100000101;end
            11'b01110010110: begin lvalue_r <= 16'b0010111100000101; rvalue_r <= 16'b0010111100010100;end
            11'b01110010111: begin lvalue_r <= 16'b0010111100010100; rvalue_r <= 16'b0010111100100010;end
            11'b01110011000: begin lvalue_r <= 16'b0010111100100010; rvalue_r <= 16'b0010111100110000;end
            11'b01110011001: begin lvalue_r <= 16'b0010111100110000; rvalue_r <= 16'b0010111100111110;end
            11'b01110011010: begin lvalue_r <= 16'b0010111100111110; rvalue_r <= 16'b0010111101001101;end
            11'b01110011011: begin lvalue_r <= 16'b0010111101001101; rvalue_r <= 16'b0010111101011011;end
            11'b01110011100: begin lvalue_r <= 16'b0010111101011011; rvalue_r <= 16'b0010111101101001;end
            11'b01110011101: begin lvalue_r <= 16'b0010111101101001; rvalue_r <= 16'b0010111101111000;end
            11'b01110011110: begin lvalue_r <= 16'b0010111101111000; rvalue_r <= 16'b0010111110000110;end
            11'b01110011111: begin lvalue_r <= 16'b0010111110000110; rvalue_r <= 16'b0010111110010100;end
            11'b01110100000: begin lvalue_r <= 16'b0010111110010100; rvalue_r <= 16'b0010111110100011;end
            11'b01110100001: begin lvalue_r <= 16'b0010111110100011; rvalue_r <= 16'b0010111110110001;end
            11'b01110100010: begin lvalue_r <= 16'b0010111110110001; rvalue_r <= 16'b0010111110111111;end
            11'b01110100011: begin lvalue_r <= 16'b0010111110111111; rvalue_r <= 16'b0010111111001101;end
            11'b01110100100: begin lvalue_r <= 16'b0010111111001101; rvalue_r <= 16'b0010111111011100;end
            11'b01110100101: begin lvalue_r <= 16'b0010111111011100; rvalue_r <= 16'b0010111111101010;end
            11'b01110100110: begin lvalue_r <= 16'b0010111111101010; rvalue_r <= 16'b0010111111111000;end
            11'b01110100111: begin lvalue_r <= 16'b0010111111111000; rvalue_r <= 16'b0011000000000111;end
            11'b01110101000: begin lvalue_r <= 16'b0011000000000111; rvalue_r <= 16'b0011000000010101;end
            11'b01110101001: begin lvalue_r <= 16'b0011000000010101; rvalue_r <= 16'b0011000000100011;end
            11'b01110101010: begin lvalue_r <= 16'b0011000000100011; rvalue_r <= 16'b0011000000110010;end
            11'b01110101011: begin lvalue_r <= 16'b0011000000110010; rvalue_r <= 16'b0011000001000000;end
            11'b01110101100: begin lvalue_r <= 16'b0011000001000000; rvalue_r <= 16'b0011000001001110;end
            11'b01110101101: begin lvalue_r <= 16'b0011000001001110; rvalue_r <= 16'b0011000001011101;end
            11'b01110101110: begin lvalue_r <= 16'b0011000001011101; rvalue_r <= 16'b0011000001101011;end
            11'b01110101111: begin lvalue_r <= 16'b0011000001101011; rvalue_r <= 16'b0011000001111010;end
            11'b01110110000: begin lvalue_r <= 16'b0011000001111010; rvalue_r <= 16'b0011000010001000;end
            11'b01110110001: begin lvalue_r <= 16'b0011000010001000; rvalue_r <= 16'b0011000010010110;end
            11'b01110110010: begin lvalue_r <= 16'b0011000010010110; rvalue_r <= 16'b0011000010100101;end
            11'b01110110011: begin lvalue_r <= 16'b0011000010100101; rvalue_r <= 16'b0011000010110011;end
            11'b01110110100: begin lvalue_r <= 16'b0011000010110011; rvalue_r <= 16'b0011000011000001;end
            11'b01110110101: begin lvalue_r <= 16'b0011000011000001; rvalue_r <= 16'b0011000011010000;end
            11'b01110110110: begin lvalue_r <= 16'b0011000011010000; rvalue_r <= 16'b0011000011011110;end
            11'b01110110111: begin lvalue_r <= 16'b0011000011011110; rvalue_r <= 16'b0011000011101101;end
            11'b01110111000: begin lvalue_r <= 16'b0011000011101101; rvalue_r <= 16'b0011000011111011;end
            11'b01110111001: begin lvalue_r <= 16'b0011000011111011; rvalue_r <= 16'b0011000100001001;end
            11'b01110111010: begin lvalue_r <= 16'b0011000100001001; rvalue_r <= 16'b0011000100011000;end
            11'b01110111011: begin lvalue_r <= 16'b0011000100011000; rvalue_r <= 16'b0011000100100110;end
            11'b01110111100: begin lvalue_r <= 16'b0011000100100110; rvalue_r <= 16'b0011000100110101;end
            11'b01110111101: begin lvalue_r <= 16'b0011000100110101; rvalue_r <= 16'b0011000101000011;end
            11'b01110111110: begin lvalue_r <= 16'b0011000101000011; rvalue_r <= 16'b0011000101010010;end
            11'b01110111111: begin lvalue_r <= 16'b0011000101010010; rvalue_r <= 16'b0011000101100000;end
            11'b01111000000: begin lvalue_r <= 16'b0011000101100000; rvalue_r <= 16'b0011000101101110;end
            11'b01111000001: begin lvalue_r <= 16'b0011000101101110; rvalue_r <= 16'b0011000101111101;end
            11'b01111000010: begin lvalue_r <= 16'b0011000101111101; rvalue_r <= 16'b0011000110001011;end
            11'b01111000011: begin lvalue_r <= 16'b0011000110001011; rvalue_r <= 16'b0011000110011010;end
            11'b01111000100: begin lvalue_r <= 16'b0011000110011010; rvalue_r <= 16'b0011000110101000;end
            11'b01111000101: begin lvalue_r <= 16'b0011000110101000; rvalue_r <= 16'b0011000110110111;end
            11'b01111000110: begin lvalue_r <= 16'b0011000110110111; rvalue_r <= 16'b0011000111000101;end
            11'b01111000111: begin lvalue_r <= 16'b0011000111000101; rvalue_r <= 16'b0011000111010100;end
            11'b01111001000: begin lvalue_r <= 16'b0011000111010100; rvalue_r <= 16'b0011000111100010;end
            11'b01111001001: begin lvalue_r <= 16'b0011000111100010; rvalue_r <= 16'b0011000111110001;end
            11'b01111001010: begin lvalue_r <= 16'b0011000111110001; rvalue_r <= 16'b0011000111111111;end
            11'b01111001011: begin lvalue_r <= 16'b0011000111111111; rvalue_r <= 16'b0011001000001110;end
            11'b01111001100: begin lvalue_r <= 16'b0011001000001110; rvalue_r <= 16'b0011001000011100;end
            11'b01111001101: begin lvalue_r <= 16'b0011001000011100; rvalue_r <= 16'b0011001000101011;end
            11'b01111001110: begin lvalue_r <= 16'b0011001000101011; rvalue_r <= 16'b0011001000111001;end
            11'b01111001111: begin lvalue_r <= 16'b0011001000111001; rvalue_r <= 16'b0011001001001000;end
            11'b01111010000: begin lvalue_r <= 16'b0011001001001000; rvalue_r <= 16'b0011001001010110;end
            11'b01111010001: begin lvalue_r <= 16'b0011001001010110; rvalue_r <= 16'b0011001001100101;end
            11'b01111010010: begin lvalue_r <= 16'b0011001001100101; rvalue_r <= 16'b0011001001110011;end
            11'b01111010011: begin lvalue_r <= 16'b0011001001110011; rvalue_r <= 16'b0011001010000010;end
            11'b01111010100: begin lvalue_r <= 16'b0011001010000010; rvalue_r <= 16'b0011001010010000;end
            11'b01111010101: begin lvalue_r <= 16'b0011001010010000; rvalue_r <= 16'b0011001010011111;end
            11'b01111010110: begin lvalue_r <= 16'b0011001010011111; rvalue_r <= 16'b0011001010101101;end
            11'b01111010111: begin lvalue_r <= 16'b0011001010101101; rvalue_r <= 16'b0011001010111100;end
            11'b01111011000: begin lvalue_r <= 16'b0011001010111100; rvalue_r <= 16'b0011001011001010;end
            11'b01111011001: begin lvalue_r <= 16'b0011001011001010; rvalue_r <= 16'b0011001011011001;end
            11'b01111011010: begin lvalue_r <= 16'b0011001011011001; rvalue_r <= 16'b0011001011100111;end
            11'b01111011011: begin lvalue_r <= 16'b0011001011100111; rvalue_r <= 16'b0011001011110110;end
            11'b01111011100: begin lvalue_r <= 16'b0011001011110110; rvalue_r <= 16'b0011001100000100;end
            11'b01111011101: begin lvalue_r <= 16'b0011001100000100; rvalue_r <= 16'b0011001100010011;end
            11'b01111011110: begin lvalue_r <= 16'b0011001100010011; rvalue_r <= 16'b0011001100100010;end
            11'b01111011111: begin lvalue_r <= 16'b0011001100100010; rvalue_r <= 16'b0011001100110000;end
            11'b01111100000: begin lvalue_r <= 16'b0011001100110000; rvalue_r <= 16'b0011001100111111;end
            11'b01111100001: begin lvalue_r <= 16'b0011001100111111; rvalue_r <= 16'b0011001101001101;end
            11'b01111100010: begin lvalue_r <= 16'b0011001101001101; rvalue_r <= 16'b0011001101011100;end
            11'b01111100011: begin lvalue_r <= 16'b0011001101011100; rvalue_r <= 16'b0011001101101011;end
            11'b01111100100: begin lvalue_r <= 16'b0011001101101011; rvalue_r <= 16'b0011001101111001;end
            11'b01111100101: begin lvalue_r <= 16'b0011001101111001; rvalue_r <= 16'b0011001110001000;end
            11'b01111100110: begin lvalue_r <= 16'b0011001110001000; rvalue_r <= 16'b0011001110010110;end
            11'b01111100111: begin lvalue_r <= 16'b0011001110010110; rvalue_r <= 16'b0011001110100101;end
            11'b01111101000: begin lvalue_r <= 16'b0011001110100101; rvalue_r <= 16'b0011001110110100;end
            11'b01111101001: begin lvalue_r <= 16'b0011001110110100; rvalue_r <= 16'b0011001111000010;end
            11'b01111101010: begin lvalue_r <= 16'b0011001111000010; rvalue_r <= 16'b0011001111010001;end
            11'b01111101011: begin lvalue_r <= 16'b0011001111010001; rvalue_r <= 16'b0011001111011111;end
            11'b01111101100: begin lvalue_r <= 16'b0011001111011111; rvalue_r <= 16'b0011001111101110;end
            11'b01111101101: begin lvalue_r <= 16'b0011001111101110; rvalue_r <= 16'b0011001111111101;end
            11'b01111101110: begin lvalue_r <= 16'b0011001111111101; rvalue_r <= 16'b0011010000001011;end
            11'b01111101111: begin lvalue_r <= 16'b0011010000001011; rvalue_r <= 16'b0011010000011010;end
            11'b01111110000: begin lvalue_r <= 16'b0011010000011010; rvalue_r <= 16'b0011010000101001;end
            11'b01111110001: begin lvalue_r <= 16'b0011010000101001; rvalue_r <= 16'b0011010000110111;end
            11'b01111110010: begin lvalue_r <= 16'b0011010000110111; rvalue_r <= 16'b0011010001000110;end
            11'b01111110011: begin lvalue_r <= 16'b0011010001000110; rvalue_r <= 16'b0011010001010101;end
            11'b01111110100: begin lvalue_r <= 16'b0011010001010101; rvalue_r <= 16'b0011010001100011;end
            11'b01111110101: begin lvalue_r <= 16'b0011010001100011; rvalue_r <= 16'b0011010001110010;end
            11'b01111110110: begin lvalue_r <= 16'b0011010001110010; rvalue_r <= 16'b0011010010000001;end
            11'b01111110111: begin lvalue_r <= 16'b0011010010000001; rvalue_r <= 16'b0011010010001111;end
            11'b01111111000: begin lvalue_r <= 16'b0011010010001111; rvalue_r <= 16'b0011010010011110;end
            11'b01111111001: begin lvalue_r <= 16'b0011010010011110; rvalue_r <= 16'b0011010010101101;end
            11'b01111111010: begin lvalue_r <= 16'b0011010010101101; rvalue_r <= 16'b0011010010111011;end
            11'b01111111011: begin lvalue_r <= 16'b0011010010111011; rvalue_r <= 16'b0011010011001010;end
            11'b01111111100: begin lvalue_r <= 16'b0011010011001010; rvalue_r <= 16'b0011010011011001;end
            11'b01111111101: begin lvalue_r <= 16'b0011010011011001; rvalue_r <= 16'b0011010011101000;end
            11'b01111111110: begin lvalue_r <= 16'b0011010011101000; rvalue_r <= 16'b0011010011110110;end
            11'b01111111111: begin lvalue_r <= 16'b0011010011110110; rvalue_r <= 16'b0011010100000101;end
            11'b10000000000: begin lvalue_r <= 16'b0011010100000101; rvalue_r <= 16'b0011010100010100;end
            11'b10000000001: begin lvalue_r <= 16'b0011010100010100; rvalue_r <= 16'b0011010100100010;end
            11'b10000000010: begin lvalue_r <= 16'b0011010100100010; rvalue_r <= 16'b0011010100110001;end
            11'b10000000011: begin lvalue_r <= 16'b0011010100110001; rvalue_r <= 16'b0011010101000000;end
            11'b10000000100: begin lvalue_r <= 16'b0011010101000000; rvalue_r <= 16'b0011010101001111;end
            11'b10000000101: begin lvalue_r <= 16'b0011010101001111; rvalue_r <= 16'b0011010101011101;end
            11'b10000000110: begin lvalue_r <= 16'b0011010101011101; rvalue_r <= 16'b0011010101101100;end
            11'b10000000111: begin lvalue_r <= 16'b0011010101101100; rvalue_r <= 16'b0011010101111011;end
            11'b10000001000: begin lvalue_r <= 16'b0011010101111011; rvalue_r <= 16'b0011010110001010;end
            11'b10000001001: begin lvalue_r <= 16'b0011010110001010; rvalue_r <= 16'b0011010110011000;end
            11'b10000001010: begin lvalue_r <= 16'b0011010110011000; rvalue_r <= 16'b0011010110100111;end
            11'b10000001011: begin lvalue_r <= 16'b0011010110100111; rvalue_r <= 16'b0011010110110110;end
            11'b10000001100: begin lvalue_r <= 16'b0011010110110110; rvalue_r <= 16'b0011010111000101;end
            11'b10000001101: begin lvalue_r <= 16'b0011010111000101; rvalue_r <= 16'b0011010111010100;end
            11'b10000001110: begin lvalue_r <= 16'b0011010111010100; rvalue_r <= 16'b0011010111100010;end
            11'b10000001111: begin lvalue_r <= 16'b0011010111100010; rvalue_r <= 16'b0011010111110001;end
            11'b10000010000: begin lvalue_r <= 16'b0011010111110001; rvalue_r <= 16'b0011011000000000;end
            11'b10000010001: begin lvalue_r <= 16'b0011011000000000; rvalue_r <= 16'b0011011000001111;end
            11'b10000010010: begin lvalue_r <= 16'b0011011000001111; rvalue_r <= 16'b0011011000011110;end
            11'b10000010011: begin lvalue_r <= 16'b0011011000011110; rvalue_r <= 16'b0011011000101100;end
            11'b10000010100: begin lvalue_r <= 16'b0011011000101100; rvalue_r <= 16'b0011011000111011;end
            11'b10000010101: begin lvalue_r <= 16'b0011011000111011; rvalue_r <= 16'b0011011001001010;end
            11'b10000010110: begin lvalue_r <= 16'b0011011001001010; rvalue_r <= 16'b0011011001011001;end
            11'b10000010111: begin lvalue_r <= 16'b0011011001011001; rvalue_r <= 16'b0011011001101000;end
            11'b10000011000: begin lvalue_r <= 16'b0011011001101000; rvalue_r <= 16'b0011011001110110;end
            11'b10000011001: begin lvalue_r <= 16'b0011011001110110; rvalue_r <= 16'b0011011010000101;end
            11'b10000011010: begin lvalue_r <= 16'b0011011010000101; rvalue_r <= 16'b0011011010010100;end
            11'b10000011011: begin lvalue_r <= 16'b0011011010010100; rvalue_r <= 16'b0011011010100011;end
            11'b10000011100: begin lvalue_r <= 16'b0011011010100011; rvalue_r <= 16'b0011011010110010;end
            11'b10000011101: begin lvalue_r <= 16'b0011011010110010; rvalue_r <= 16'b0011011011000001;end
            11'b10000011110: begin lvalue_r <= 16'b0011011011000001; rvalue_r <= 16'b0011011011010000;end
            11'b10000011111: begin lvalue_r <= 16'b0011011011010000; rvalue_r <= 16'b0011011011011110;end
            11'b10000100000: begin lvalue_r <= 16'b0011011011011110; rvalue_r <= 16'b0011011011101101;end
            11'b10000100001: begin lvalue_r <= 16'b0011011011101101; rvalue_r <= 16'b0011011011111100;end
            11'b10000100010: begin lvalue_r <= 16'b0011011011111100; rvalue_r <= 16'b0011011100001011;end
            11'b10000100011: begin lvalue_r <= 16'b0011011100001011; rvalue_r <= 16'b0011011100011010;end
            11'b10000100100: begin lvalue_r <= 16'b0011011100011010; rvalue_r <= 16'b0011011100101001;end
            11'b10000100101: begin lvalue_r <= 16'b0011011100101001; rvalue_r <= 16'b0011011100111000;end
            11'b10000100110: begin lvalue_r <= 16'b0011011100111000; rvalue_r <= 16'b0011011101000111;end
            11'b10000100111: begin lvalue_r <= 16'b0011011101000111; rvalue_r <= 16'b0011011101010110;end
            11'b10000101000: begin lvalue_r <= 16'b0011011101010110; rvalue_r <= 16'b0011011101100101;end
            11'b10000101001: begin lvalue_r <= 16'b0011011101100101; rvalue_r <= 16'b0011011101110011;end
            11'b10000101010: begin lvalue_r <= 16'b0011011101110011; rvalue_r <= 16'b0011011110000010;end
            11'b10000101011: begin lvalue_r <= 16'b0011011110000010; rvalue_r <= 16'b0011011110010001;end
            11'b10000101100: begin lvalue_r <= 16'b0011011110010001; rvalue_r <= 16'b0011011110100000;end
            11'b10000101101: begin lvalue_r <= 16'b0011011110100000; rvalue_r <= 16'b0011011110101111;end
            11'b10000101110: begin lvalue_r <= 16'b0011011110101111; rvalue_r <= 16'b0011011110111110;end
            11'b10000101111: begin lvalue_r <= 16'b0011011110111110; rvalue_r <= 16'b0011011111001101;end
            11'b10000110000: begin lvalue_r <= 16'b0011011111001101; rvalue_r <= 16'b0011011111011100;end
            11'b10000110001: begin lvalue_r <= 16'b0011011111011100; rvalue_r <= 16'b0011011111101011;end
            11'b10000110010: begin lvalue_r <= 16'b0011011111101011; rvalue_r <= 16'b0011011111111010;end
            11'b10000110011: begin lvalue_r <= 16'b0011011111111010; rvalue_r <= 16'b0011100000001001;end
            11'b10000110100: begin lvalue_r <= 16'b0011100000001001; rvalue_r <= 16'b0011100000011000;end
            11'b10000110101: begin lvalue_r <= 16'b0011100000011000; rvalue_r <= 16'b0011100000100111;end
            11'b10000110110: begin lvalue_r <= 16'b0011100000100111; rvalue_r <= 16'b0011100000110110;end
            11'b10000110111: begin lvalue_r <= 16'b0011100000110110; rvalue_r <= 16'b0011100001000101;end
            11'b10000111000: begin lvalue_r <= 16'b0011100001000101; rvalue_r <= 16'b0011100001010100;end
            11'b10000111001: begin lvalue_r <= 16'b0011100001010100; rvalue_r <= 16'b0011100001100011;end
            11'b10000111010: begin lvalue_r <= 16'b0011100001100011; rvalue_r <= 16'b0011100001110010;end
            11'b10000111011: begin lvalue_r <= 16'b0011100001110010; rvalue_r <= 16'b0011100010000001;end
            11'b10000111100: begin lvalue_r <= 16'b0011100010000001; rvalue_r <= 16'b0011100010010000;end
            11'b10000111101: begin lvalue_r <= 16'b0011100010010000; rvalue_r <= 16'b0011100010011111;end
            11'b10000111110: begin lvalue_r <= 16'b0011100010011111; rvalue_r <= 16'b0011100010101110;end
            11'b10000111111: begin lvalue_r <= 16'b0011100010101110; rvalue_r <= 16'b0011100010111101;end
            11'b10001000000: begin lvalue_r <= 16'b0011100010111101; rvalue_r <= 16'b0011100011001100;end
            11'b10001000001: begin lvalue_r <= 16'b0011100011001100; rvalue_r <= 16'b0011100011011011;end
            11'b10001000010: begin lvalue_r <= 16'b0011100011011011; rvalue_r <= 16'b0011100011101010;end
            11'b10001000011: begin lvalue_r <= 16'b0011100011101010; rvalue_r <= 16'b0011100011111001;end
            11'b10001000100: begin lvalue_r <= 16'b0011100011111001; rvalue_r <= 16'b0011100100001000;end
            11'b10001000101: begin lvalue_r <= 16'b0011100100001000; rvalue_r <= 16'b0011100100010111;end
            11'b10001000110: begin lvalue_r <= 16'b0011100100010111; rvalue_r <= 16'b0011100100100110;end
            11'b10001000111: begin lvalue_r <= 16'b0011100100100110; rvalue_r <= 16'b0011100100110110;end
            11'b10001001000: begin lvalue_r <= 16'b0011100100110110; rvalue_r <= 16'b0011100101000101;end
            11'b10001001001: begin lvalue_r <= 16'b0011100101000101; rvalue_r <= 16'b0011100101010100;end
            11'b10001001010: begin lvalue_r <= 16'b0011100101010100; rvalue_r <= 16'b0011100101100011;end
            11'b10001001011: begin lvalue_r <= 16'b0011100101100011; rvalue_r <= 16'b0011100101110010;end
            11'b10001001100: begin lvalue_r <= 16'b0011100101110010; rvalue_r <= 16'b0011100110000001;end
            11'b10001001101: begin lvalue_r <= 16'b0011100110000001; rvalue_r <= 16'b0011100110010000;end
            11'b10001001110: begin lvalue_r <= 16'b0011100110010000; rvalue_r <= 16'b0011100110011111;end
            11'b10001001111: begin lvalue_r <= 16'b0011100110011111; rvalue_r <= 16'b0011100110101110;end
            11'b10001010000: begin lvalue_r <= 16'b0011100110101110; rvalue_r <= 16'b0011100110111101;end
            11'b10001010001: begin lvalue_r <= 16'b0011100110111101; rvalue_r <= 16'b0011100111001101;end
            11'b10001010010: begin lvalue_r <= 16'b0011100111001101; rvalue_r <= 16'b0011100111011100;end
            11'b10001010011: begin lvalue_r <= 16'b0011100111011100; rvalue_r <= 16'b0011100111101011;end
            11'b10001010100: begin lvalue_r <= 16'b0011100111101011; rvalue_r <= 16'b0011100111111010;end
            11'b10001010101: begin lvalue_r <= 16'b0011100111111010; rvalue_r <= 16'b0011101000001001;end
            11'b10001010110: begin lvalue_r <= 16'b0011101000001001; rvalue_r <= 16'b0011101000011000;end
            11'b10001010111: begin lvalue_r <= 16'b0011101000011000; rvalue_r <= 16'b0011101000100111;end
            11'b10001011000: begin lvalue_r <= 16'b0011101000100111; rvalue_r <= 16'b0011101000110111;end
            11'b10001011001: begin lvalue_r <= 16'b0011101000110111; rvalue_r <= 16'b0011101001000110;end
            11'b10001011010: begin lvalue_r <= 16'b0011101001000110; rvalue_r <= 16'b0011101001010101;end
            11'b10001011011: begin lvalue_r <= 16'b0011101001010101; rvalue_r <= 16'b0011101001100100;end
            11'b10001011100: begin lvalue_r <= 16'b0011101001100100; rvalue_r <= 16'b0011101001110011;end
            11'b10001011101: begin lvalue_r <= 16'b0011101001110011; rvalue_r <= 16'b0011101010000010;end
            11'b10001011110: begin lvalue_r <= 16'b0011101010000010; rvalue_r <= 16'b0011101010010010;end
            11'b10001011111: begin lvalue_r <= 16'b0011101010010010; rvalue_r <= 16'b0011101010100001;end
            11'b10001100000: begin lvalue_r <= 16'b0011101010100001; rvalue_r <= 16'b0011101010110000;end
            11'b10001100001: begin lvalue_r <= 16'b0011101010110000; rvalue_r <= 16'b0011101010111111;end
            11'b10001100010: begin lvalue_r <= 16'b0011101010111111; rvalue_r <= 16'b0011101011001110;end
            11'b10001100011: begin lvalue_r <= 16'b0011101011001110; rvalue_r <= 16'b0011101011011110;end
            11'b10001100100: begin lvalue_r <= 16'b0011101011011110; rvalue_r <= 16'b0011101011101101;end
            11'b10001100101: begin lvalue_r <= 16'b0011101011101101; rvalue_r <= 16'b0011101011111100;end
            11'b10001100110: begin lvalue_r <= 16'b0011101011111100; rvalue_r <= 16'b0011101100001011;end
            11'b10001100111: begin lvalue_r <= 16'b0011101100001011; rvalue_r <= 16'b0011101100011011;end
            11'b10001101000: begin lvalue_r <= 16'b0011101100011011; rvalue_r <= 16'b0011101100101010;end
            11'b10001101001: begin lvalue_r <= 16'b0011101100101010; rvalue_r <= 16'b0011101100111001;end
            11'b10001101010: begin lvalue_r <= 16'b0011101100111001; rvalue_r <= 16'b0011101101001000;end
            11'b10001101011: begin lvalue_r <= 16'b0011101101001000; rvalue_r <= 16'b0011101101011000;end
            11'b10001101100: begin lvalue_r <= 16'b0011101101011000; rvalue_r <= 16'b0011101101100111;end
            11'b10001101101: begin lvalue_r <= 16'b0011101101100111; rvalue_r <= 16'b0011101101110110;end
            11'b10001101110: begin lvalue_r <= 16'b0011101101110110; rvalue_r <= 16'b0011101110000101;end
            11'b10001101111: begin lvalue_r <= 16'b0011101110000101; rvalue_r <= 16'b0011101110010101;end
            11'b10001110000: begin lvalue_r <= 16'b0011101110010101; rvalue_r <= 16'b0011101110100100;end
            11'b10001110001: begin lvalue_r <= 16'b0011101110100100; rvalue_r <= 16'b0011101110110011;end
            11'b10001110010: begin lvalue_r <= 16'b0011101110110011; rvalue_r <= 16'b0011101111000011;end
            11'b10001110011: begin lvalue_r <= 16'b0011101111000011; rvalue_r <= 16'b0011101111010010;end
            11'b10001110100: begin lvalue_r <= 16'b0011101111010010; rvalue_r <= 16'b0011101111100001;end
            11'b10001110101: begin lvalue_r <= 16'b0011101111100001; rvalue_r <= 16'b0011101111110001;end
            11'b10001110110: begin lvalue_r <= 16'b0011101111110001; rvalue_r <= 16'b0011110000000000;end
            11'b10001110111: begin lvalue_r <= 16'b0011110000000000; rvalue_r <= 16'b0011110000001111;end
            11'b10001111000: begin lvalue_r <= 16'b0011110000001111; rvalue_r <= 16'b0011110000011111;end
            11'b10001111001: begin lvalue_r <= 16'b0011110000011111; rvalue_r <= 16'b0011110000101110;end
            11'b10001111010: begin lvalue_r <= 16'b0011110000101110; rvalue_r <= 16'b0011110000111101;end
            11'b10001111011: begin lvalue_r <= 16'b0011110000111101; rvalue_r <= 16'b0011110001001101;end
            11'b10001111100: begin lvalue_r <= 16'b0011110001001101; rvalue_r <= 16'b0011110001011100;end
            11'b10001111101: begin lvalue_r <= 16'b0011110001011100; rvalue_r <= 16'b0011110001101011;end
            11'b10001111110: begin lvalue_r <= 16'b0011110001101011; rvalue_r <= 16'b0011110001111011;end
            11'b10001111111: begin lvalue_r <= 16'b0011110001111011; rvalue_r <= 16'b0011110010001010;end
            11'b10010000000: begin lvalue_r <= 16'b0011110010001010; rvalue_r <= 16'b0011110010011001;end
            11'b10010000001: begin lvalue_r <= 16'b0011110010011001; rvalue_r <= 16'b0011110010101001;end
            11'b10010000010: begin lvalue_r <= 16'b0011110010101001; rvalue_r <= 16'b0011110010111000;end
            11'b10010000011: begin lvalue_r <= 16'b0011110010111000; rvalue_r <= 16'b0011110011001000;end
            11'b10010000100: begin lvalue_r <= 16'b0011110011001000; rvalue_r <= 16'b0011110011010111;end
            11'b10010000101: begin lvalue_r <= 16'b0011110011010111; rvalue_r <= 16'b0011110011100110;end
            11'b10010000110: begin lvalue_r <= 16'b0011110011100110; rvalue_r <= 16'b0011110011110110;end
            11'b10010000111: begin lvalue_r <= 16'b0011110011110110; rvalue_r <= 16'b0011110100000101;end
            11'b10010001000: begin lvalue_r <= 16'b0011110100000101; rvalue_r <= 16'b0011110100010101;end
            11'b10010001001: begin lvalue_r <= 16'b0011110100010101; rvalue_r <= 16'b0011110100100100;end
            11'b10010001010: begin lvalue_r <= 16'b0011110100100100; rvalue_r <= 16'b0011110100110100;end
            11'b10010001011: begin lvalue_r <= 16'b0011110100110100; rvalue_r <= 16'b0011110101000011;end
            11'b10010001100: begin lvalue_r <= 16'b0011110101000011; rvalue_r <= 16'b0011110101010010;end
            11'b10010001101: begin lvalue_r <= 16'b0011110101010010; rvalue_r <= 16'b0011110101100010;end
            11'b10010001110: begin lvalue_r <= 16'b0011110101100010; rvalue_r <= 16'b0011110101110001;end
            11'b10010001111: begin lvalue_r <= 16'b0011110101110001; rvalue_r <= 16'b0011110110000001;end
            11'b10010010000: begin lvalue_r <= 16'b0011110110000001; rvalue_r <= 16'b0011110110010000;end
            11'b10010010001: begin lvalue_r <= 16'b0011110110010000; rvalue_r <= 16'b0011110110100000;end
            11'b10010010010: begin lvalue_r <= 16'b0011110110100000; rvalue_r <= 16'b0011110110101111;end
            11'b10010010011: begin lvalue_r <= 16'b0011110110101111; rvalue_r <= 16'b0011110110111111;end
            11'b10010010100: begin lvalue_r <= 16'b0011110110111111; rvalue_r <= 16'b0011110111001110;end
            11'b10010010101: begin lvalue_r <= 16'b0011110111001110; rvalue_r <= 16'b0011110111011110;end
            11'b10010010110: begin lvalue_r <= 16'b0011110111011110; rvalue_r <= 16'b0011110111101101;end
            11'b10010010111: begin lvalue_r <= 16'b0011110111101101; rvalue_r <= 16'b0011110111111101;end
            11'b10010011000: begin lvalue_r <= 16'b0011110111111101; rvalue_r <= 16'b0011111000001100;end
            11'b10010011001: begin lvalue_r <= 16'b0011111000001100; rvalue_r <= 16'b0011111000011100;end
            11'b10010011010: begin lvalue_r <= 16'b0011111000011100; rvalue_r <= 16'b0011111000101011;end
            11'b10010011011: begin lvalue_r <= 16'b0011111000101011; rvalue_r <= 16'b0011111000111011;end
            11'b10010011100: begin lvalue_r <= 16'b0011111000111011; rvalue_r <= 16'b0011111001001010;end
            11'b10010011101: begin lvalue_r <= 16'b0011111001001010; rvalue_r <= 16'b0011111001011010;end
            11'b10010011110: begin lvalue_r <= 16'b0011111001011010; rvalue_r <= 16'b0011111001101010;end
            11'b10010011111: begin lvalue_r <= 16'b0011111001101010; rvalue_r <= 16'b0011111001111001;end
            11'b10010100000: begin lvalue_r <= 16'b0011111001111001; rvalue_r <= 16'b0011111010001001;end
            11'b10010100001: begin lvalue_r <= 16'b0011111010001001; rvalue_r <= 16'b0011111010011000;end
            11'b10010100010: begin lvalue_r <= 16'b0011111010011000; rvalue_r <= 16'b0011111010101000;end
            11'b10010100011: begin lvalue_r <= 16'b0011111010101000; rvalue_r <= 16'b0011111010110111;end
            11'b10010100100: begin lvalue_r <= 16'b0011111010110111; rvalue_r <= 16'b0011111011000111;end
            11'b10010100101: begin lvalue_r <= 16'b0011111011000111; rvalue_r <= 16'b0011111011010111;end
            11'b10010100110: begin lvalue_r <= 16'b0011111011010111; rvalue_r <= 16'b0011111011100110;end
            11'b10010100111: begin lvalue_r <= 16'b0011111011100110; rvalue_r <= 16'b0011111011110110;end
            11'b10010101000: begin lvalue_r <= 16'b0011111011110110; rvalue_r <= 16'b0011111100000101;end
            11'b10010101001: begin lvalue_r <= 16'b0011111100000101; rvalue_r <= 16'b0011111100010101;end
            11'b10010101010: begin lvalue_r <= 16'b0011111100010101; rvalue_r <= 16'b0011111100100101;end
            11'b10010101011: begin lvalue_r <= 16'b0011111100100101; rvalue_r <= 16'b0011111100110100;end
            11'b10010101100: begin lvalue_r <= 16'b0011111100110100; rvalue_r <= 16'b0011111101000100;end
            11'b10010101101: begin lvalue_r <= 16'b0011111101000100; rvalue_r <= 16'b0011111101010011;end
            11'b10010101110: begin lvalue_r <= 16'b0011111101010011; rvalue_r <= 16'b0011111101100011;end
            11'b10010101111: begin lvalue_r <= 16'b0011111101100011; rvalue_r <= 16'b0011111101110011;end
            11'b10010110000: begin lvalue_r <= 16'b0011111101110011; rvalue_r <= 16'b0011111110000010;end
            11'b10010110001: begin lvalue_r <= 16'b0011111110000010; rvalue_r <= 16'b0011111110010010;end
            11'b10010110010: begin lvalue_r <= 16'b0011111110010010; rvalue_r <= 16'b0011111110100010;end
            11'b10010110011: begin lvalue_r <= 16'b0011111110100010; rvalue_r <= 16'b0011111110110001;end
            11'b10010110100: begin lvalue_r <= 16'b0011111110110001; rvalue_r <= 16'b0011111111000001;end
            11'b10010110101: begin lvalue_r <= 16'b0011111111000001; rvalue_r <= 16'b0011111111010001;end
            11'b10010110110: begin lvalue_r <= 16'b0011111111010001; rvalue_r <= 16'b0011111111100001;end
            11'b10010110111: begin lvalue_r <= 16'b0011111111100001; rvalue_r <= 16'b0011111111110000;end
            11'b10010111000: begin lvalue_r <= 16'b0011111111110000; rvalue_r <= 16'b0100000000000000;end
            11'b10010111001: begin lvalue_r <= 16'b0100000000000000; rvalue_r <= 16'b0100000000010000;end
            11'b10010111010: begin lvalue_r <= 16'b0100000000010000; rvalue_r <= 16'b0100000000011111;end
            11'b10010111011: begin lvalue_r <= 16'b0100000000011111; rvalue_r <= 16'b0100000000101111;end
            11'b10010111100: begin lvalue_r <= 16'b0100000000101111; rvalue_r <= 16'b0100000000111111;end
            11'b10010111101: begin lvalue_r <= 16'b0100000000111111; rvalue_r <= 16'b0100000001001111;end
            11'b10010111110: begin lvalue_r <= 16'b0100000001001111; rvalue_r <= 16'b0100000001011110;end
            11'b10010111111: begin lvalue_r <= 16'b0100000001011110; rvalue_r <= 16'b0100000001101110;end
            11'b10011000000: begin lvalue_r <= 16'b0100000001101110; rvalue_r <= 16'b0100000001111110;end
            11'b10011000001: begin lvalue_r <= 16'b0100000001111110; rvalue_r <= 16'b0100000010001110;end
            11'b10011000010: begin lvalue_r <= 16'b0100000010001110; rvalue_r <= 16'b0100000010011101;end
            11'b10011000011: begin lvalue_r <= 16'b0100000010011101; rvalue_r <= 16'b0100000010101101;end
            11'b10011000100: begin lvalue_r <= 16'b0100000010101101; rvalue_r <= 16'b0100000010111101;end
            11'b10011000101: begin lvalue_r <= 16'b0100000010111101; rvalue_r <= 16'b0100000011001101;end
            11'b10011000110: begin lvalue_r <= 16'b0100000011001101; rvalue_r <= 16'b0100000011011100;end
            11'b10011000111: begin lvalue_r <= 16'b0100000011011100; rvalue_r <= 16'b0100000011101100;end
            11'b10011001000: begin lvalue_r <= 16'b0100000011101100; rvalue_r <= 16'b0100000011111100;end
            11'b10011001001: begin lvalue_r <= 16'b0100000011111100; rvalue_r <= 16'b0100000100001100;end
            11'b10011001010: begin lvalue_r <= 16'b0100000100001100; rvalue_r <= 16'b0100000100011100;end
            11'b10011001011: begin lvalue_r <= 16'b0100000100011100; rvalue_r <= 16'b0100000100101011;end
            11'b10011001100: begin lvalue_r <= 16'b0100000100101011; rvalue_r <= 16'b0100000100111011;end
            11'b10011001101: begin lvalue_r <= 16'b0100000100111011; rvalue_r <= 16'b0100000101001011;end
            11'b10011001110: begin lvalue_r <= 16'b0100000101001011; rvalue_r <= 16'b0100000101011011;end
            11'b10011001111: begin lvalue_r <= 16'b0100000101011011; rvalue_r <= 16'b0100000101101011;end
            11'b10011010000: begin lvalue_r <= 16'b0100000101101011; rvalue_r <= 16'b0100000101111011;end
            11'b10011010001: begin lvalue_r <= 16'b0100000101111011; rvalue_r <= 16'b0100000110001011;end
            11'b10011010010: begin lvalue_r <= 16'b0100000110001011; rvalue_r <= 16'b0100000110011010;end
            11'b10011010011: begin lvalue_r <= 16'b0100000110011010; rvalue_r <= 16'b0100000110101010;end
            11'b10011010100: begin lvalue_r <= 16'b0100000110101010; rvalue_r <= 16'b0100000110111010;end
            11'b10011010101: begin lvalue_r <= 16'b0100000110111010; rvalue_r <= 16'b0100000111001010;end
            11'b10011010110: begin lvalue_r <= 16'b0100000111001010; rvalue_r <= 16'b0100000111011010;end
            11'b10011010111: begin lvalue_r <= 16'b0100000111011010; rvalue_r <= 16'b0100000111101010;end
            11'b10011011000: begin lvalue_r <= 16'b0100000111101010; rvalue_r <= 16'b0100000111111010;end
            11'b10011011001: begin lvalue_r <= 16'b0100000111111010; rvalue_r <= 16'b0100001000001010;end
            11'b10011011010: begin lvalue_r <= 16'b0100001000001010; rvalue_r <= 16'b0100001000011010;end
            11'b10011011011: begin lvalue_r <= 16'b0100001000011010; rvalue_r <= 16'b0100001000101001;end
            11'b10011011100: begin lvalue_r <= 16'b0100001000101001; rvalue_r <= 16'b0100001000111001;end
            11'b10011011101: begin lvalue_r <= 16'b0100001000111001; rvalue_r <= 16'b0100001001001001;end
            11'b10011011110: begin lvalue_r <= 16'b0100001001001001; rvalue_r <= 16'b0100001001011001;end
            11'b10011011111: begin lvalue_r <= 16'b0100001001011001; rvalue_r <= 16'b0100001001101001;end
            11'b10011100000: begin lvalue_r <= 16'b0100001001101001; rvalue_r <= 16'b0100001001111001;end
            11'b10011100001: begin lvalue_r <= 16'b0100001001111001; rvalue_r <= 16'b0100001010001001;end
            11'b10011100010: begin lvalue_r <= 16'b0100001010001001; rvalue_r <= 16'b0100001010011001;end
            11'b10011100011: begin lvalue_r <= 16'b0100001010011001; rvalue_r <= 16'b0100001010101001;end
            11'b10011100100: begin lvalue_r <= 16'b0100001010101001; rvalue_r <= 16'b0100001010111001;end
            11'b10011100101: begin lvalue_r <= 16'b0100001010111001; rvalue_r <= 16'b0100001011001001;end
            11'b10011100110: begin lvalue_r <= 16'b0100001011001001; rvalue_r <= 16'b0100001011011001;end
            11'b10011100111: begin lvalue_r <= 16'b0100001011011001; rvalue_r <= 16'b0100001011101001;end
            11'b10011101000: begin lvalue_r <= 16'b0100001011101001; rvalue_r <= 16'b0100001011111001;end
            11'b10011101001: begin lvalue_r <= 16'b0100001011111001; rvalue_r <= 16'b0100001100001001;end
            11'b10011101010: begin lvalue_r <= 16'b0100001100001001; rvalue_r <= 16'b0100001100011001;end
            11'b10011101011: begin lvalue_r <= 16'b0100001100011001; rvalue_r <= 16'b0100001100101001;end
            11'b10011101100: begin lvalue_r <= 16'b0100001100101001; rvalue_r <= 16'b0100001100111001;end
            11'b10011101101: begin lvalue_r <= 16'b0100001100111001; rvalue_r <= 16'b0100001101001001;end
            11'b10011101110: begin lvalue_r <= 16'b0100001101001001; rvalue_r <= 16'b0100001101011001;end
            11'b10011101111: begin lvalue_r <= 16'b0100001101011001; rvalue_r <= 16'b0100001101101001;end
            11'b10011110000: begin lvalue_r <= 16'b0100001101101001; rvalue_r <= 16'b0100001101111001;end
            11'b10011110001: begin lvalue_r <= 16'b0100001101111001; rvalue_r <= 16'b0100001110001001;end
            11'b10011110010: begin lvalue_r <= 16'b0100001110001001; rvalue_r <= 16'b0100001110011001;end
            11'b10011110011: begin lvalue_r <= 16'b0100001110011001; rvalue_r <= 16'b0100001110101001;end
            11'b10011110100: begin lvalue_r <= 16'b0100001110101001; rvalue_r <= 16'b0100001110111010;end
            11'b10011110101: begin lvalue_r <= 16'b0100001110111010; rvalue_r <= 16'b0100001111001010;end
            11'b10011110110: begin lvalue_r <= 16'b0100001111001010; rvalue_r <= 16'b0100001111011010;end
            11'b10011110111: begin lvalue_r <= 16'b0100001111011010; rvalue_r <= 16'b0100001111101010;end
            11'b10011111000: begin lvalue_r <= 16'b0100001111101010; rvalue_r <= 16'b0100001111111010;end
            11'b10011111001: begin lvalue_r <= 16'b0100001111111010; rvalue_r <= 16'b0100010000001010;end
            11'b10011111010: begin lvalue_r <= 16'b0100010000001010; rvalue_r <= 16'b0100010000011010;end
            11'b10011111011: begin lvalue_r <= 16'b0100010000011010; rvalue_r <= 16'b0100010000101010;end
            11'b10011111100: begin lvalue_r <= 16'b0100010000101010; rvalue_r <= 16'b0100010000111010;end
            11'b10011111101: begin lvalue_r <= 16'b0100010000111010; rvalue_r <= 16'b0100010001001011;end
            11'b10011111110: begin lvalue_r <= 16'b0100010001001011; rvalue_r <= 16'b0100010001011011;end
            11'b10011111111: begin lvalue_r <= 16'b0100010001011011; rvalue_r <= 16'b0100010001101011;end
            11'b10100000000: begin lvalue_r <= 16'b0100010001101011; rvalue_r <= 16'b0100010001111011;end
            11'b10100000001: begin lvalue_r <= 16'b0100010001111011; rvalue_r <= 16'b0100010010001011;end
            11'b10100000010: begin lvalue_r <= 16'b0100010010001011; rvalue_r <= 16'b0100010010011011;end
            11'b10100000011: begin lvalue_r <= 16'b0100010010011011; rvalue_r <= 16'b0100010010101100;end
            11'b10100000100: begin lvalue_r <= 16'b0100010010101100; rvalue_r <= 16'b0100010010111100;end
            11'b10100000101: begin lvalue_r <= 16'b0100010010111100; rvalue_r <= 16'b0100010011001100;end
            11'b10100000110: begin lvalue_r <= 16'b0100010011001100; rvalue_r <= 16'b0100010011011100;end
            11'b10100000111: begin lvalue_r <= 16'b0100010011011100; rvalue_r <= 16'b0100010011101100;end
            11'b10100001000: begin lvalue_r <= 16'b0100010011101100; rvalue_r <= 16'b0100010011111101;end
            11'b10100001001: begin lvalue_r <= 16'b0100010011111101; rvalue_r <= 16'b0100010100001101;end
            11'b10100001010: begin lvalue_r <= 16'b0100010100001101; rvalue_r <= 16'b0100010100011101;end
            11'b10100001011: begin lvalue_r <= 16'b0100010100011101; rvalue_r <= 16'b0100010100101101;end
            11'b10100001100: begin lvalue_r <= 16'b0100010100101101; rvalue_r <= 16'b0100010100111101;end
            11'b10100001101: begin lvalue_r <= 16'b0100010100111101; rvalue_r <= 16'b0100010101001110;end
            11'b10100001110: begin lvalue_r <= 16'b0100010101001110; rvalue_r <= 16'b0100010101011110;end
            11'b10100001111: begin lvalue_r <= 16'b0100010101011110; rvalue_r <= 16'b0100010101101110;end
            11'b10100010000: begin lvalue_r <= 16'b0100010101101110; rvalue_r <= 16'b0100010101111110;end
            11'b10100010001: begin lvalue_r <= 16'b0100010101111110; rvalue_r <= 16'b0100010110001111;end
            11'b10100010010: begin lvalue_r <= 16'b0100010110001111; rvalue_r <= 16'b0100010110011111;end
            11'b10100010011: begin lvalue_r <= 16'b0100010110011111; rvalue_r <= 16'b0100010110101111;end
            11'b10100010100: begin lvalue_r <= 16'b0100010110101111; rvalue_r <= 16'b0100010111000000;end
            11'b10100010101: begin lvalue_r <= 16'b0100010111000000; rvalue_r <= 16'b0100010111010000;end
            11'b10100010110: begin lvalue_r <= 16'b0100010111010000; rvalue_r <= 16'b0100010111100000;end
            11'b10100010111: begin lvalue_r <= 16'b0100010111100000; rvalue_r <= 16'b0100010111110001;end
            11'b10100011000: begin lvalue_r <= 16'b0100010111110001; rvalue_r <= 16'b0100011000000001;end
            11'b10100011001: begin lvalue_r <= 16'b0100011000000001; rvalue_r <= 16'b0100011000010001;end
            11'b10100011010: begin lvalue_r <= 16'b0100011000010001; rvalue_r <= 16'b0100011000100010;end
            11'b10100011011: begin lvalue_r <= 16'b0100011000100010; rvalue_r <= 16'b0100011000110010;end
            11'b10100011100: begin lvalue_r <= 16'b0100011000110010; rvalue_r <= 16'b0100011001000010;end
            11'b10100011101: begin lvalue_r <= 16'b0100011001000010; rvalue_r <= 16'b0100011001010011;end
            11'b10100011110: begin lvalue_r <= 16'b0100011001010011; rvalue_r <= 16'b0100011001100011;end
            11'b10100011111: begin lvalue_r <= 16'b0100011001100011; rvalue_r <= 16'b0100011001110011;end
            11'b10100100000: begin lvalue_r <= 16'b0100011001110011; rvalue_r <= 16'b0100011010000100;end
            11'b10100100001: begin lvalue_r <= 16'b0100011010000100; rvalue_r <= 16'b0100011010010100;end
            11'b10100100010: begin lvalue_r <= 16'b0100011010010100; rvalue_r <= 16'b0100011010100100;end
            11'b10100100011: begin lvalue_r <= 16'b0100011010100100; rvalue_r <= 16'b0100011010110101;end
            11'b10100100100: begin lvalue_r <= 16'b0100011010110101; rvalue_r <= 16'b0100011011000101;end
            11'b10100100101: begin lvalue_r <= 16'b0100011011000101; rvalue_r <= 16'b0100011011010110;end
            11'b10100100110: begin lvalue_r <= 16'b0100011011010110; rvalue_r <= 16'b0100011011100110;end
            11'b10100100111: begin lvalue_r <= 16'b0100011011100110; rvalue_r <= 16'b0100011011110111;end
            11'b10100101000: begin lvalue_r <= 16'b0100011011110111; rvalue_r <= 16'b0100011100000111;end
            11'b10100101001: begin lvalue_r <= 16'b0100011100000111; rvalue_r <= 16'b0100011100010111;end
            11'b10100101010: begin lvalue_r <= 16'b0100011100010111; rvalue_r <= 16'b0100011100101000;end
            11'b10100101011: begin lvalue_r <= 16'b0100011100101000; rvalue_r <= 16'b0100011100111000;end
            11'b10100101100: begin lvalue_r <= 16'b0100011100111000; rvalue_r <= 16'b0100011101001001;end
            11'b10100101101: begin lvalue_r <= 16'b0100011101001001; rvalue_r <= 16'b0100011101011001;end
            11'b10100101110: begin lvalue_r <= 16'b0100011101011001; rvalue_r <= 16'b0100011101101010;end
            11'b10100101111: begin lvalue_r <= 16'b0100011101101010; rvalue_r <= 16'b0100011101111010;end
            11'b10100110000: begin lvalue_r <= 16'b0100011101111010; rvalue_r <= 16'b0100011110001011;end
            11'b10100110001: begin lvalue_r <= 16'b0100011110001011; rvalue_r <= 16'b0100011110011011;end
            11'b10100110010: begin lvalue_r <= 16'b0100011110011011; rvalue_r <= 16'b0100011110101100;end
            11'b10100110011: begin lvalue_r <= 16'b0100011110101100; rvalue_r <= 16'b0100011110111100;end
            11'b10100110100: begin lvalue_r <= 16'b0100011110111100; rvalue_r <= 16'b0100011111001101;end
            11'b10100110101: begin lvalue_r <= 16'b0100011111001101; rvalue_r <= 16'b0100011111011101;end
            11'b10100110110: begin lvalue_r <= 16'b0100011111011101; rvalue_r <= 16'b0100011111101110;end
            11'b10100110111: begin lvalue_r <= 16'b0100011111101110; rvalue_r <= 16'b0100011111111110;end
            11'b10100111000: begin lvalue_r <= 16'b0100011111111110; rvalue_r <= 16'b0100100000001111;end
            11'b10100111001: begin lvalue_r <= 16'b0100100000001111; rvalue_r <= 16'b0100100000011111;end
            11'b10100111010: begin lvalue_r <= 16'b0100100000011111; rvalue_r <= 16'b0100100000110000;end
            11'b10100111011: begin lvalue_r <= 16'b0100100000110000; rvalue_r <= 16'b0100100001000001;end
            11'b10100111100: begin lvalue_r <= 16'b0100100001000001; rvalue_r <= 16'b0100100001010001;end
            11'b10100111101: begin lvalue_r <= 16'b0100100001010001; rvalue_r <= 16'b0100100001100010;end
            11'b10100111110: begin lvalue_r <= 16'b0100100001100010; rvalue_r <= 16'b0100100001110010;end
            11'b10100111111: begin lvalue_r <= 16'b0100100001110010; rvalue_r <= 16'b0100100010000011;end
            11'b10101000000: begin lvalue_r <= 16'b0100100010000011; rvalue_r <= 16'b0100100010010011;end
            11'b10101000001: begin lvalue_r <= 16'b0100100010010011; rvalue_r <= 16'b0100100010100100;end
            11'b10101000010: begin lvalue_r <= 16'b0100100010100100; rvalue_r <= 16'b0100100010110101;end
            11'b10101000011: begin lvalue_r <= 16'b0100100010110101; rvalue_r <= 16'b0100100011000101;end
            11'b10101000100: begin lvalue_r <= 16'b0100100011000101; rvalue_r <= 16'b0100100011010110;end
            11'b10101000101: begin lvalue_r <= 16'b0100100011010110; rvalue_r <= 16'b0100100011100111;end
            11'b10101000110: begin lvalue_r <= 16'b0100100011100111; rvalue_r <= 16'b0100100011110111;end
            11'b10101000111: begin lvalue_r <= 16'b0100100011110111; rvalue_r <= 16'b0100100100001000;end
            11'b10101001000: begin lvalue_r <= 16'b0100100100001000; rvalue_r <= 16'b0100100100011001;end
            11'b10101001001: begin lvalue_r <= 16'b0100100100011001; rvalue_r <= 16'b0100100100101001;end
            11'b10101001010: begin lvalue_r <= 16'b0100100100101001; rvalue_r <= 16'b0100100100111010;end
            11'b10101001011: begin lvalue_r <= 16'b0100100100111010; rvalue_r <= 16'b0100100101001011;end
            11'b10101001100: begin lvalue_r <= 16'b0100100101001011; rvalue_r <= 16'b0100100101011011;end
            11'b10101001101: begin lvalue_r <= 16'b0100100101011011; rvalue_r <= 16'b0100100101101100;end
            11'b10101001110: begin lvalue_r <= 16'b0100100101101100; rvalue_r <= 16'b0100100101111101;end
            11'b10101001111: begin lvalue_r <= 16'b0100100101111101; rvalue_r <= 16'b0100100110001101;end
            11'b10101010000: begin lvalue_r <= 16'b0100100110001101; rvalue_r <= 16'b0100100110011110;end
            11'b10101010001: begin lvalue_r <= 16'b0100100110011110; rvalue_r <= 16'b0100100110101111;end
            11'b10101010010: begin lvalue_r <= 16'b0100100110101111; rvalue_r <= 16'b0100100111000000;end
            11'b10101010011: begin lvalue_r <= 16'b0100100111000000; rvalue_r <= 16'b0100100111010000;end
            11'b10101010100: begin lvalue_r <= 16'b0100100111010000; rvalue_r <= 16'b0100100111100001;end
            11'b10101010101: begin lvalue_r <= 16'b0100100111100001; rvalue_r <= 16'b0100100111110010;end
            11'b10101010110: begin lvalue_r <= 16'b0100100111110010; rvalue_r <= 16'b0100101000000011;end
            11'b10101010111: begin lvalue_r <= 16'b0100101000000011; rvalue_r <= 16'b0100101000010011;end
            11'b10101011000: begin lvalue_r <= 16'b0100101000010011; rvalue_r <= 16'b0100101000100100;end
            11'b10101011001: begin lvalue_r <= 16'b0100101000100100; rvalue_r <= 16'b0100101000110101;end
            11'b10101011010: begin lvalue_r <= 16'b0100101000110101; rvalue_r <= 16'b0100101001000110;end
            11'b10101011011: begin lvalue_r <= 16'b0100101001000110; rvalue_r <= 16'b0100101001010110;end
            11'b10101011100: begin lvalue_r <= 16'b0100101001010110; rvalue_r <= 16'b0100101001100111;end
            11'b10101011101: begin lvalue_r <= 16'b0100101001100111; rvalue_r <= 16'b0100101001111000;end
            11'b10101011110: begin lvalue_r <= 16'b0100101001111000; rvalue_r <= 16'b0100101010001001;end
            11'b10101011111: begin lvalue_r <= 16'b0100101010001001; rvalue_r <= 16'b0100101010011010;end
            11'b10101100000: begin lvalue_r <= 16'b0100101010011010; rvalue_r <= 16'b0100101010101011;end
            11'b10101100001: begin lvalue_r <= 16'b0100101010101011; rvalue_r <= 16'b0100101010111011;end
            11'b10101100010: begin lvalue_r <= 16'b0100101010111011; rvalue_r <= 16'b0100101011001100;end
            11'b10101100011: begin lvalue_r <= 16'b0100101011001100; rvalue_r <= 16'b0100101011011101;end
            11'b10101100100: begin lvalue_r <= 16'b0100101011011101; rvalue_r <= 16'b0100101011101110;end
            11'b10101100101: begin lvalue_r <= 16'b0100101011101110; rvalue_r <= 16'b0100101011111111;end
            11'b10101100110: begin lvalue_r <= 16'b0100101011111111; rvalue_r <= 16'b0100101100010000;end
            11'b10101100111: begin lvalue_r <= 16'b0100101100010000; rvalue_r <= 16'b0100101100100001;end
            11'b10101101000: begin lvalue_r <= 16'b0100101100100001; rvalue_r <= 16'b0100101100110010;end
            11'b10101101001: begin lvalue_r <= 16'b0100101100110010; rvalue_r <= 16'b0100101101000010;end
            11'b10101101010: begin lvalue_r <= 16'b0100101101000010; rvalue_r <= 16'b0100101101010011;end
            11'b10101101011: begin lvalue_r <= 16'b0100101101010011; rvalue_r <= 16'b0100101101100100;end
            11'b10101101100: begin lvalue_r <= 16'b0100101101100100; rvalue_r <= 16'b0100101101110101;end
            11'b10101101101: begin lvalue_r <= 16'b0100101101110101; rvalue_r <= 16'b0100101110000110;end
            11'b10101101110: begin lvalue_r <= 16'b0100101110000110; rvalue_r <= 16'b0100101110010111;end
            11'b10101101111: begin lvalue_r <= 16'b0100101110010111; rvalue_r <= 16'b0100101110101000;end
            11'b10101110000: begin lvalue_r <= 16'b0100101110101000; rvalue_r <= 16'b0100101110111001;end
            11'b10101110001: begin lvalue_r <= 16'b0100101110111001; rvalue_r <= 16'b0100101111001010;end
            11'b10101110010: begin lvalue_r <= 16'b0100101111001010; rvalue_r <= 16'b0100101111011011;end
            11'b10101110011: begin lvalue_r <= 16'b0100101111011011; rvalue_r <= 16'b0100101111101100;end
            11'b10101110100: begin lvalue_r <= 16'b0100101111101100; rvalue_r <= 16'b0100101111111101;end
            11'b10101110101: begin lvalue_r <= 16'b0100101111111101; rvalue_r <= 16'b0100110000001110;end
            11'b10101110110: begin lvalue_r <= 16'b0100110000001110; rvalue_r <= 16'b0100110000011111;end
            11'b10101110111: begin lvalue_r <= 16'b0100110000011111; rvalue_r <= 16'b0100110000110000;end
            11'b10101111000: begin lvalue_r <= 16'b0100110000110000; rvalue_r <= 16'b0100110001000001;end
            11'b10101111001: begin lvalue_r <= 16'b0100110001000001; rvalue_r <= 16'b0100110001010010;end
            11'b10101111010: begin lvalue_r <= 16'b0100110001010010; rvalue_r <= 16'b0100110001100011;end
            11'b10101111011: begin lvalue_r <= 16'b0100110001100011; rvalue_r <= 16'b0100110001110100;end
            11'b10101111100: begin lvalue_r <= 16'b0100110001110100; rvalue_r <= 16'b0100110010000101;end
            11'b10101111101: begin lvalue_r <= 16'b0100110010000101; rvalue_r <= 16'b0100110010010110;end
            11'b10101111110: begin lvalue_r <= 16'b0100110010010110; rvalue_r <= 16'b0100110010100111;end
            11'b10101111111: begin lvalue_r <= 16'b0100110010100111; rvalue_r <= 16'b0100110010111000;end
            11'b10110000000: begin lvalue_r <= 16'b0100110010111000; rvalue_r <= 16'b0100110011001001;end
            11'b10110000001: begin lvalue_r <= 16'b0100110011001001; rvalue_r <= 16'b0100110011011011;end
            11'b10110000010: begin lvalue_r <= 16'b0100110011011011; rvalue_r <= 16'b0100110011101100;end
            11'b10110000011: begin lvalue_r <= 16'b0100110011101100; rvalue_r <= 16'b0100110011111101;end
            11'b10110000100: begin lvalue_r <= 16'b0100110011111101; rvalue_r <= 16'b0100110100001110;end
            11'b10110000101: begin lvalue_r <= 16'b0100110100001110; rvalue_r <= 16'b0100110100011111;end
            11'b10110000110: begin lvalue_r <= 16'b0100110100011111; rvalue_r <= 16'b0100110100110000;end
            11'b10110000111: begin lvalue_r <= 16'b0100110100110000; rvalue_r <= 16'b0100110101000001;end
            11'b10110001000: begin lvalue_r <= 16'b0100110101000001; rvalue_r <= 16'b0100110101010010;end
            11'b10110001001: begin lvalue_r <= 16'b0100110101010010; rvalue_r <= 16'b0100110101100100;end
            11'b10110001010: begin lvalue_r <= 16'b0100110101100100; rvalue_r <= 16'b0100110101110101;end
            11'b10110001011: begin lvalue_r <= 16'b0100110101110101; rvalue_r <= 16'b0100110110000110;end
            11'b10110001100: begin lvalue_r <= 16'b0100110110000110; rvalue_r <= 16'b0100110110010111;end
            11'b10110001101: begin lvalue_r <= 16'b0100110110010111; rvalue_r <= 16'b0100110110101000;end
            11'b10110001110: begin lvalue_r <= 16'b0100110110101000; rvalue_r <= 16'b0100110110111001;end
            11'b10110001111: begin lvalue_r <= 16'b0100110110111001; rvalue_r <= 16'b0100110111001011;end
            11'b10110010000: begin lvalue_r <= 16'b0100110111001011; rvalue_r <= 16'b0100110111011100;end
            11'b10110010001: begin lvalue_r <= 16'b0100110111011100; rvalue_r <= 16'b0100110111101101;end
            11'b10110010010: begin lvalue_r <= 16'b0100110111101101; rvalue_r <= 16'b0100110111111110;end
            11'b10110010011: begin lvalue_r <= 16'b0100110111111110; rvalue_r <= 16'b0100111000010000;end
            11'b10110010100: begin lvalue_r <= 16'b0100111000010000; rvalue_r <= 16'b0100111000100001;end
            11'b10110010101: begin lvalue_r <= 16'b0100111000100001; rvalue_r <= 16'b0100111000110010;end
            11'b10110010110: begin lvalue_r <= 16'b0100111000110010; rvalue_r <= 16'b0100111001000011;end
            11'b10110010111: begin lvalue_r <= 16'b0100111001000011; rvalue_r <= 16'b0100111001010101;end
            11'b10110011000: begin lvalue_r <= 16'b0100111001010101; rvalue_r <= 16'b0100111001100110;end
            11'b10110011001: begin lvalue_r <= 16'b0100111001100110; rvalue_r <= 16'b0100111001110111;end
            11'b10110011010: begin lvalue_r <= 16'b0100111001110111; rvalue_r <= 16'b0100111010001000;end
            11'b10110011011: begin lvalue_r <= 16'b0100111010001000; rvalue_r <= 16'b0100111010011010;end
            11'b10110011100: begin lvalue_r <= 16'b0100111010011010; rvalue_r <= 16'b0100111010101011;end
            11'b10110011101: begin lvalue_r <= 16'b0100111010101011; rvalue_r <= 16'b0100111010111100;end
            11'b10110011110: begin lvalue_r <= 16'b0100111010111100; rvalue_r <= 16'b0100111011001110;end
            11'b10110011111: begin lvalue_r <= 16'b0100111011001110; rvalue_r <= 16'b0100111011011111;end
            11'b10110100000: begin lvalue_r <= 16'b0100111011011111; rvalue_r <= 16'b0100111011110000;end
            11'b10110100001: begin lvalue_r <= 16'b0100111011110000; rvalue_r <= 16'b0100111100000010;end
            11'b10110100010: begin lvalue_r <= 16'b0100111100000010; rvalue_r <= 16'b0100111100010011;end
            11'b10110100011: begin lvalue_r <= 16'b0100111100010011; rvalue_r <= 16'b0100111100100100;end
            11'b10110100100: begin lvalue_r <= 16'b0100111100100100; rvalue_r <= 16'b0100111100110110;end
            11'b10110100101: begin lvalue_r <= 16'b0100111100110110; rvalue_r <= 16'b0100111101000111;end
            11'b10110100110: begin lvalue_r <= 16'b0100111101000111; rvalue_r <= 16'b0100111101011001;end
            11'b10110100111: begin lvalue_r <= 16'b0100111101011001; rvalue_r <= 16'b0100111101101010;end
            11'b10110101000: begin lvalue_r <= 16'b0100111101101010; rvalue_r <= 16'b0100111101111011;end
            11'b10110101001: begin lvalue_r <= 16'b0100111101111011; rvalue_r <= 16'b0100111110001101;end
            11'b10110101010: begin lvalue_r <= 16'b0100111110001101; rvalue_r <= 16'b0100111110011110;end
            11'b10110101011: begin lvalue_r <= 16'b0100111110011110; rvalue_r <= 16'b0100111110110000;end
            11'b10110101100: begin lvalue_r <= 16'b0100111110110000; rvalue_r <= 16'b0100111111000001;end
            11'b10110101101: begin lvalue_r <= 16'b0100111111000001; rvalue_r <= 16'b0100111111010011;end
            11'b10110101110: begin lvalue_r <= 16'b0100111111010011; rvalue_r <= 16'b0100111111100100;end
            11'b10110101111: begin lvalue_r <= 16'b0100111111100100; rvalue_r <= 16'b0100111111110110;end
            11'b10110110000: begin lvalue_r <= 16'b0100111111110110; rvalue_r <= 16'b0101000000000111;end
            11'b10110110001: begin lvalue_r <= 16'b0101000000000111; rvalue_r <= 16'b0101000000011000;end
            11'b10110110010: begin lvalue_r <= 16'b0101000000011000; rvalue_r <= 16'b0101000000101010;end
            11'b10110110011: begin lvalue_r <= 16'b0101000000101010; rvalue_r <= 16'b0101000000111011;end
            11'b10110110100: begin lvalue_r <= 16'b0101000000111011; rvalue_r <= 16'b0101000001001101;end
            11'b10110110101: begin lvalue_r <= 16'b0101000001001101; rvalue_r <= 16'b0101000001011110;end
            11'b10110110110: begin lvalue_r <= 16'b0101000001011110; rvalue_r <= 16'b0101000001110000;end
            11'b10110110111: begin lvalue_r <= 16'b0101000001110000; rvalue_r <= 16'b0101000010000010;end
            11'b10110111000: begin lvalue_r <= 16'b0101000010000010; rvalue_r <= 16'b0101000010010011;end
            11'b10110111001: begin lvalue_r <= 16'b0101000010010011; rvalue_r <= 16'b0101000010100101;end
            11'b10110111010: begin lvalue_r <= 16'b0101000010100101; rvalue_r <= 16'b0101000010110110;end
            11'b10110111011: begin lvalue_r <= 16'b0101000010110110; rvalue_r <= 16'b0101000011001000;end
            11'b10110111100: begin lvalue_r <= 16'b0101000011001000; rvalue_r <= 16'b0101000011011001;end
            11'b10110111101: begin lvalue_r <= 16'b0101000011011001; rvalue_r <= 16'b0101000011101011;end
            11'b10110111110: begin lvalue_r <= 16'b0101000011101011; rvalue_r <= 16'b0101000011111101;end
            11'b10110111111: begin lvalue_r <= 16'b0101000011111101; rvalue_r <= 16'b0101000100001110;end
            11'b10111000000: begin lvalue_r <= 16'b0101000100001110; rvalue_r <= 16'b0101000100100000;end
            11'b10111000001: begin lvalue_r <= 16'b0101000100100000; rvalue_r <= 16'b0101000100110001;end
            11'b10111000010: begin lvalue_r <= 16'b0101000100110001; rvalue_r <= 16'b0101000101000011;end
            11'b10111000011: begin lvalue_r <= 16'b0101000101000011; rvalue_r <= 16'b0101000101010101;end
            11'b10111000100: begin lvalue_r <= 16'b0101000101010101; rvalue_r <= 16'b0101000101100110;end
            11'b10111000101: begin lvalue_r <= 16'b0101000101100110; rvalue_r <= 16'b0101000101111000;end
            11'b10111000110: begin lvalue_r <= 16'b0101000101111000; rvalue_r <= 16'b0101000110001010;end
            11'b10111000111: begin lvalue_r <= 16'b0101000110001010; rvalue_r <= 16'b0101000110011011;end
            11'b10111001000: begin lvalue_r <= 16'b0101000110011011; rvalue_r <= 16'b0101000110101101;end
            11'b10111001001: begin lvalue_r <= 16'b0101000110101101; rvalue_r <= 16'b0101000110111111;end
            11'b10111001010: begin lvalue_r <= 16'b0101000110111111; rvalue_r <= 16'b0101000111010000;end
            11'b10111001011: begin lvalue_r <= 16'b0101000111010000; rvalue_r <= 16'b0101000111100010;end
            11'b10111001100: begin lvalue_r <= 16'b0101000111100010; rvalue_r <= 16'b0101000111110100;end
            11'b10111001101: begin lvalue_r <= 16'b0101000111110100; rvalue_r <= 16'b0101001000000101;end
            11'b10111001110: begin lvalue_r <= 16'b0101001000000101; rvalue_r <= 16'b0101001000010111;end
            11'b10111001111: begin lvalue_r <= 16'b0101001000010111; rvalue_r <= 16'b0101001000101001;end
            11'b10111010000: begin lvalue_r <= 16'b0101001000101001; rvalue_r <= 16'b0101001000111011;end
            11'b10111010001: begin lvalue_r <= 16'b0101001000111011; rvalue_r <= 16'b0101001001001100;end
            11'b10111010010: begin lvalue_r <= 16'b0101001001001100; rvalue_r <= 16'b0101001001011110;end
            11'b10111010011: begin lvalue_r <= 16'b0101001001011110; rvalue_r <= 16'b0101001001110000;end
            11'b10111010100: begin lvalue_r <= 16'b0101001001110000; rvalue_r <= 16'b0101001010000010;end
            11'b10111010101: begin lvalue_r <= 16'b0101001010000010; rvalue_r <= 16'b0101001010010100;end
            11'b10111010110: begin lvalue_r <= 16'b0101001010010100; rvalue_r <= 16'b0101001010100101;end
            11'b10111010111: begin lvalue_r <= 16'b0101001010100101; rvalue_r <= 16'b0101001010110111;end
            11'b10111011000: begin lvalue_r <= 16'b0101001010110111; rvalue_r <= 16'b0101001011001001;end
            11'b10111011001: begin lvalue_r <= 16'b0101001011001001; rvalue_r <= 16'b0101001011011011;end
            11'b10111011010: begin lvalue_r <= 16'b0101001011011011; rvalue_r <= 16'b0101001011101101;end
            11'b10111011011: begin lvalue_r <= 16'b0101001011101101; rvalue_r <= 16'b0101001011111110;end
            11'b10111011100: begin lvalue_r <= 16'b0101001011111110; rvalue_r <= 16'b0101001100010000;end
            11'b10111011101: begin lvalue_r <= 16'b0101001100010000; rvalue_r <= 16'b0101001100100010;end
            11'b10111011110: begin lvalue_r <= 16'b0101001100100010; rvalue_r <= 16'b0101001100110100;end
            11'b10111011111: begin lvalue_r <= 16'b0101001100110100; rvalue_r <= 16'b0101001101000110;end
            11'b10111100000: begin lvalue_r <= 16'b0101001101000110; rvalue_r <= 16'b0101001101011000;end
            11'b10111100001: begin lvalue_r <= 16'b0101001101011000; rvalue_r <= 16'b0101001101101010;end
            11'b10111100010: begin lvalue_r <= 16'b0101001101101010; rvalue_r <= 16'b0101001101111100;end
            11'b10111100011: begin lvalue_r <= 16'b0101001101111100; rvalue_r <= 16'b0101001110001110;end
            11'b10111100100: begin lvalue_r <= 16'b0101001110001110; rvalue_r <= 16'b0101001110011111;end
            11'b10111100101: begin lvalue_r <= 16'b0101001110011111; rvalue_r <= 16'b0101001110110001;end
            11'b10111100110: begin lvalue_r <= 16'b0101001110110001; rvalue_r <= 16'b0101001111000011;end
            11'b10111100111: begin lvalue_r <= 16'b0101001111000011; rvalue_r <= 16'b0101001111010101;end
            11'b10111101000: begin lvalue_r <= 16'b0101001111010101; rvalue_r <= 16'b0101001111100111;end
            11'b10111101001: begin lvalue_r <= 16'b0101001111100111; rvalue_r <= 16'b0101001111111001;end
            11'b10111101010: begin lvalue_r <= 16'b0101001111111001; rvalue_r <= 16'b0101010000001011;end
            11'b10111101011: begin lvalue_r <= 16'b0101010000001011; rvalue_r <= 16'b0101010000011101;end
            11'b10111101100: begin lvalue_r <= 16'b0101010000011101; rvalue_r <= 16'b0101010000101111;end
            11'b10111101101: begin lvalue_r <= 16'b0101010000101111; rvalue_r <= 16'b0101010001000001;end
            11'b10111101110: begin lvalue_r <= 16'b0101010001000001; rvalue_r <= 16'b0101010001010011;end
            11'b10111101111: begin lvalue_r <= 16'b0101010001010011; rvalue_r <= 16'b0101010001100101;end
            11'b10111110000: begin lvalue_r <= 16'b0101010001100101; rvalue_r <= 16'b0101010001110111;end
            11'b10111110001: begin lvalue_r <= 16'b0101010001110111; rvalue_r <= 16'b0101010010001001;end
            11'b10111110010: begin lvalue_r <= 16'b0101010010001001; rvalue_r <= 16'b0101010010011011;end
            11'b10111110011: begin lvalue_r <= 16'b0101010010011011; rvalue_r <= 16'b0101010010101101;end
            11'b10111110100: begin lvalue_r <= 16'b0101010010101101; rvalue_r <= 16'b0101010010111111;end
            11'b10111110101: begin lvalue_r <= 16'b0101010010111111; rvalue_r <= 16'b0101010011010010;end
            11'b10111110110: begin lvalue_r <= 16'b0101010011010010; rvalue_r <= 16'b0101010011100100;end
            11'b10111110111: begin lvalue_r <= 16'b0101010011100100; rvalue_r <= 16'b0101010011110110;end
            11'b10111111000: begin lvalue_r <= 16'b0101010011110110; rvalue_r <= 16'b0101010100001000;end
            11'b10111111001: begin lvalue_r <= 16'b0101010100001000; rvalue_r <= 16'b0101010100011010;end
            11'b10111111010: begin lvalue_r <= 16'b0101010100011010; rvalue_r <= 16'b0101010100101100;end
            11'b10111111011: begin lvalue_r <= 16'b0101010100101100; rvalue_r <= 16'b0101010100111110;end
            11'b10111111100: begin lvalue_r <= 16'b0101010100111110; rvalue_r <= 16'b0101010101010000;end
            11'b10111111101: begin lvalue_r <= 16'b0101010101010000; rvalue_r <= 16'b0101010101100011;end
            11'b10111111110: begin lvalue_r <= 16'b0101010101100011; rvalue_r <= 16'b0101010101110101;end
            11'b10111111111: begin lvalue_r <= 16'b0101010101110101; rvalue_r <= 16'b0101010110000111;end
            11'b11000000000: begin lvalue_r <= 16'b0101010110000111; rvalue_r <= 16'b0101010110011001;end
            11'b11000000001: begin lvalue_r <= 16'b0101010110011001; rvalue_r <= 16'b0101010110101011;end
            11'b11000000010: begin lvalue_r <= 16'b0101010110101011; rvalue_r <= 16'b0101010110111101;end
            11'b11000000011: begin lvalue_r <= 16'b0101010110111101; rvalue_r <= 16'b0101010111010000;end
            11'b11000000100: begin lvalue_r <= 16'b0101010111010000; rvalue_r <= 16'b0101010111100010;end
            11'b11000000101: begin lvalue_r <= 16'b0101010111100010; rvalue_r <= 16'b0101010111110100;end
            11'b11000000110: begin lvalue_r <= 16'b0101010111110100; rvalue_r <= 16'b0101011000000110;end
            11'b11000000111: begin lvalue_r <= 16'b0101011000000110; rvalue_r <= 16'b0101011000011001;end
            11'b11000001000: begin lvalue_r <= 16'b0101011000011001; rvalue_r <= 16'b0101011000101011;end
            11'b11000001001: begin lvalue_r <= 16'b0101011000101011; rvalue_r <= 16'b0101011000111101;end
            11'b11000001010: begin lvalue_r <= 16'b0101011000111101; rvalue_r <= 16'b0101011001001111;end
            11'b11000001011: begin lvalue_r <= 16'b0101011001001111; rvalue_r <= 16'b0101011001100010;end
            11'b11000001100: begin lvalue_r <= 16'b0101011001100010; rvalue_r <= 16'b0101011001110100;end
            11'b11000001101: begin lvalue_r <= 16'b0101011001110100; rvalue_r <= 16'b0101011010000110;end
            11'b11000001110: begin lvalue_r <= 16'b0101011010000110; rvalue_r <= 16'b0101011010011001;end
            11'b11000001111: begin lvalue_r <= 16'b0101011010011001; rvalue_r <= 16'b0101011010101011;end
            11'b11000010000: begin lvalue_r <= 16'b0101011010101011; rvalue_r <= 16'b0101011010111101;end
            11'b11000010001: begin lvalue_r <= 16'b0101011010111101; rvalue_r <= 16'b0101011011010000;end
            11'b11000010010: begin lvalue_r <= 16'b0101011011010000; rvalue_r <= 16'b0101011011100010;end
            11'b11000010011: begin lvalue_r <= 16'b0101011011100010; rvalue_r <= 16'b0101011011110100;end
            11'b11000010100: begin lvalue_r <= 16'b0101011011110100; rvalue_r <= 16'b0101011100000111;end
            11'b11000010101: begin lvalue_r <= 16'b0101011100000111; rvalue_r <= 16'b0101011100011001;end
            11'b11000010110: begin lvalue_r <= 16'b0101011100011001; rvalue_r <= 16'b0101011100101011;end
            11'b11000010111: begin lvalue_r <= 16'b0101011100101011; rvalue_r <= 16'b0101011100111110;end
            11'b11000011000: begin lvalue_r <= 16'b0101011100111110; rvalue_r <= 16'b0101011101010000;end
            11'b11000011001: begin lvalue_r <= 16'b0101011101010000; rvalue_r <= 16'b0101011101100011;end
            11'b11000011010: begin lvalue_r <= 16'b0101011101100011; rvalue_r <= 16'b0101011101110101;end
            11'b11000011011: begin lvalue_r <= 16'b0101011101110101; rvalue_r <= 16'b0101011110001000;end
            11'b11000011100: begin lvalue_r <= 16'b0101011110001000; rvalue_r <= 16'b0101011110011010;end
            11'b11000011101: begin lvalue_r <= 16'b0101011110011010; rvalue_r <= 16'b0101011110101100;end
            11'b11000011110: begin lvalue_r <= 16'b0101011110101100; rvalue_r <= 16'b0101011110111111;end
            11'b11000011111: begin lvalue_r <= 16'b0101011110111111; rvalue_r <= 16'b0101011111010001;end
            11'b11000100000: begin lvalue_r <= 16'b0101011111010001; rvalue_r <= 16'b0101011111100100;end
            11'b11000100001: begin lvalue_r <= 16'b0101011111100100; rvalue_r <= 16'b0101011111110110;end
            11'b11000100010: begin lvalue_r <= 16'b0101011111110110; rvalue_r <= 16'b0101100000001001;end
            11'b11000100011: begin lvalue_r <= 16'b0101100000001001; rvalue_r <= 16'b0101100000011011;end
            11'b11000100100: begin lvalue_r <= 16'b0101100000011011; rvalue_r <= 16'b0101100000101110;end
            11'b11000100101: begin lvalue_r <= 16'b0101100000101110; rvalue_r <= 16'b0101100001000000;end
            11'b11000100110: begin lvalue_r <= 16'b0101100001000000; rvalue_r <= 16'b0101100001010011;end
            11'b11000100111: begin lvalue_r <= 16'b0101100001010011; rvalue_r <= 16'b0101100001100110;end
            11'b11000101000: begin lvalue_r <= 16'b0101100001100110; rvalue_r <= 16'b0101100001111000;end
            11'b11000101001: begin lvalue_r <= 16'b0101100001111000; rvalue_r <= 16'b0101100010001011;end
            11'b11000101010: begin lvalue_r <= 16'b0101100010001011; rvalue_r <= 16'b0101100010011101;end
            11'b11000101011: begin lvalue_r <= 16'b0101100010011101; rvalue_r <= 16'b0101100010110000;end
            11'b11000101100: begin lvalue_r <= 16'b0101100010110000; rvalue_r <= 16'b0101100011000010;end
            11'b11000101101: begin lvalue_r <= 16'b0101100011000010; rvalue_r <= 16'b0101100011010101;end
            11'b11000101110: begin lvalue_r <= 16'b0101100011010101; rvalue_r <= 16'b0101100011101000;end
            11'b11000101111: begin lvalue_r <= 16'b0101100011101000; rvalue_r <= 16'b0101100011111010;end
            11'b11000110000: begin lvalue_r <= 16'b0101100011111010; rvalue_r <= 16'b0101100100001101;end
            11'b11000110001: begin lvalue_r <= 16'b0101100100001101; rvalue_r <= 16'b0101100100100000;end
            11'b11000110010: begin lvalue_r <= 16'b0101100100100000; rvalue_r <= 16'b0101100100110010;end
            11'b11000110011: begin lvalue_r <= 16'b0101100100110010; rvalue_r <= 16'b0101100101000101;end
            11'b11000110100: begin lvalue_r <= 16'b0101100101000101; rvalue_r <= 16'b0101100101011000;end
            11'b11000110101: begin lvalue_r <= 16'b0101100101011000; rvalue_r <= 16'b0101100101101010;end
            11'b11000110110: begin lvalue_r <= 16'b0101100101101010; rvalue_r <= 16'b0101100101111101;end
            11'b11000110111: begin lvalue_r <= 16'b0101100101111101; rvalue_r <= 16'b0101100110010000;end
            11'b11000111000: begin lvalue_r <= 16'b0101100110010000; rvalue_r <= 16'b0101100110100010;end
            11'b11000111001: begin lvalue_r <= 16'b0101100110100010; rvalue_r <= 16'b0101100110110101;end
            11'b11000111010: begin lvalue_r <= 16'b0101100110110101; rvalue_r <= 16'b0101100111001000;end
            11'b11000111011: begin lvalue_r <= 16'b0101100111001000; rvalue_r <= 16'b0101100111011011;end
            11'b11000111100: begin lvalue_r <= 16'b0101100111011011; rvalue_r <= 16'b0101100111101101;end
            11'b11000111101: begin lvalue_r <= 16'b0101100111101101; rvalue_r <= 16'b0101101000000000;end
            11'b11000111110: begin lvalue_r <= 16'b0101101000000000; rvalue_r <= 16'b0101101000010011;end
            11'b11000111111: begin lvalue_r <= 16'b0101101000010011; rvalue_r <= 16'b0101101000100110;end
            11'b11001000000: begin lvalue_r <= 16'b0101101000100110; rvalue_r <= 16'b0101101000111001;end
            11'b11001000001: begin lvalue_r <= 16'b0101101000111001; rvalue_r <= 16'b0101101001001011;end
            11'b11001000010: begin lvalue_r <= 16'b0101101001001011; rvalue_r <= 16'b0101101001011110;end
            11'b11001000011: begin lvalue_r <= 16'b0101101001011110; rvalue_r <= 16'b0101101001110001;end
            11'b11001000100: begin lvalue_r <= 16'b0101101001110001; rvalue_r <= 16'b0101101010000100;end
            11'b11001000101: begin lvalue_r <= 16'b0101101010000100; rvalue_r <= 16'b0101101010010111;end
            11'b11001000110: begin lvalue_r <= 16'b0101101010010111; rvalue_r <= 16'b0101101010101010;end
            11'b11001000111: begin lvalue_r <= 16'b0101101010101010; rvalue_r <= 16'b0101101010111101;end
            11'b11001001000: begin lvalue_r <= 16'b0101101010111101; rvalue_r <= 16'b0101101011001111;end
            11'b11001001001: begin lvalue_r <= 16'b0101101011001111; rvalue_r <= 16'b0101101011100010;end
            11'b11001001010: begin lvalue_r <= 16'b0101101011100010; rvalue_r <= 16'b0101101011110101;end
            11'b11001001011: begin lvalue_r <= 16'b0101101011110101; rvalue_r <= 16'b0101101100001000;end
            11'b11001001100: begin lvalue_r <= 16'b0101101100001000; rvalue_r <= 16'b0101101100011011;end
            11'b11001001101: begin lvalue_r <= 16'b0101101100011011; rvalue_r <= 16'b0101101100101110;end
            11'b11001001110: begin lvalue_r <= 16'b0101101100101110; rvalue_r <= 16'b0101101101000001;end
            11'b11001001111: begin lvalue_r <= 16'b0101101101000001; rvalue_r <= 16'b0101101101010100;end
            11'b11001010000: begin lvalue_r <= 16'b0101101101010100; rvalue_r <= 16'b0101101101100111;end
            11'b11001010001: begin lvalue_r <= 16'b0101101101100111; rvalue_r <= 16'b0101101101111010;end
            11'b11001010010: begin lvalue_r <= 16'b0101101101111010; rvalue_r <= 16'b0101101110001101;end
            11'b11001010011: begin lvalue_r <= 16'b0101101110001101; rvalue_r <= 16'b0101101110100000;end
            11'b11001010100: begin lvalue_r <= 16'b0101101110100000; rvalue_r <= 16'b0101101110110011;end
            11'b11001010101: begin lvalue_r <= 16'b0101101110110011; rvalue_r <= 16'b0101101111000110;end
            11'b11001010110: begin lvalue_r <= 16'b0101101111000110; rvalue_r <= 16'b0101101111011001;end
            11'b11001010111: begin lvalue_r <= 16'b0101101111011001; rvalue_r <= 16'b0101101111101100;end
            11'b11001011000: begin lvalue_r <= 16'b0101101111101100; rvalue_r <= 16'b0101101111111111;end
            11'b11001011001: begin lvalue_r <= 16'b0101101111111111; rvalue_r <= 16'b0101110000010010;end
            11'b11001011010: begin lvalue_r <= 16'b0101110000010010; rvalue_r <= 16'b0101110000100101;end
            11'b11001011011: begin lvalue_r <= 16'b0101110000100101; rvalue_r <= 16'b0101110000111000;end
            11'b11001011100: begin lvalue_r <= 16'b0101110000111000; rvalue_r <= 16'b0101110001001011;end
            11'b11001011101: begin lvalue_r <= 16'b0101110001001011; rvalue_r <= 16'b0101110001011110;end
            11'b11001011110: begin lvalue_r <= 16'b0101110001011110; rvalue_r <= 16'b0101110001110010;end
            11'b11001011111: begin lvalue_r <= 16'b0101110001110010; rvalue_r <= 16'b0101110010000101;end
            11'b11001100000: begin lvalue_r <= 16'b0101110010000101; rvalue_r <= 16'b0101110010011000;end
            11'b11001100001: begin lvalue_r <= 16'b0101110010011000; rvalue_r <= 16'b0101110010101011;end
            11'b11001100010: begin lvalue_r <= 16'b0101110010101011; rvalue_r <= 16'b0101110010111110;end
            11'b11001100011: begin lvalue_r <= 16'b0101110010111110; rvalue_r <= 16'b0101110011010001;end
            11'b11001100100: begin lvalue_r <= 16'b0101110011010001; rvalue_r <= 16'b0101110011100100;end
            11'b11001100101: begin lvalue_r <= 16'b0101110011100100; rvalue_r <= 16'b0101110011111000;end
            11'b11001100110: begin lvalue_r <= 16'b0101110011111000; rvalue_r <= 16'b0101110100001011;end
            11'b11001100111: begin lvalue_r <= 16'b0101110100001011; rvalue_r <= 16'b0101110100011110;end
            11'b11001101000: begin lvalue_r <= 16'b0101110100011110; rvalue_r <= 16'b0101110100110001;end
            11'b11001101001: begin lvalue_r <= 16'b0101110100110001; rvalue_r <= 16'b0101110101000101;end
            11'b11001101010: begin lvalue_r <= 16'b0101110101000101; rvalue_r <= 16'b0101110101011000;end
            11'b11001101011: begin lvalue_r <= 16'b0101110101011000; rvalue_r <= 16'b0101110101101011;end
            11'b11001101100: begin lvalue_r <= 16'b0101110101101011; rvalue_r <= 16'b0101110101111110;end
            11'b11001101101: begin lvalue_r <= 16'b0101110101111110; rvalue_r <= 16'b0101110110010010;end
            11'b11001101110: begin lvalue_r <= 16'b0101110110010010; rvalue_r <= 16'b0101110110100101;end
            11'b11001101111: begin lvalue_r <= 16'b0101110110100101; rvalue_r <= 16'b0101110110111000;end
            11'b11001110000: begin lvalue_r <= 16'b0101110110111000; rvalue_r <= 16'b0101110111001011;end
            11'b11001110001: begin lvalue_r <= 16'b0101110111001011; rvalue_r <= 16'b0101110111011111;end
            11'b11001110010: begin lvalue_r <= 16'b0101110111011111; rvalue_r <= 16'b0101110111110010;end
            11'b11001110011: begin lvalue_r <= 16'b0101110111110010; rvalue_r <= 16'b0101111000000101;end
            11'b11001110100: begin lvalue_r <= 16'b0101111000000101; rvalue_r <= 16'b0101111000011001;end
            11'b11001110101: begin lvalue_r <= 16'b0101111000011001; rvalue_r <= 16'b0101111000101100;end
            11'b11001110110: begin lvalue_r <= 16'b0101111000101100; rvalue_r <= 16'b0101111001000000;end
            11'b11001110111: begin lvalue_r <= 16'b0101111001000000; rvalue_r <= 16'b0101111001010011;end
            11'b11001111000: begin lvalue_r <= 16'b0101111001010011; rvalue_r <= 16'b0101111001100110;end
            11'b11001111001: begin lvalue_r <= 16'b0101111001100110; rvalue_r <= 16'b0101111001111010;end
            11'b11001111010: begin lvalue_r <= 16'b0101111001111010; rvalue_r <= 16'b0101111010001101;end
            11'b11001111011: begin lvalue_r <= 16'b0101111010001101; rvalue_r <= 16'b0101111010100001;end
            11'b11001111100: begin lvalue_r <= 16'b0101111010100001; rvalue_r <= 16'b0101111010110100;end
            11'b11001111101: begin lvalue_r <= 16'b0101111010110100; rvalue_r <= 16'b0101111011000111;end
            11'b11001111110: begin lvalue_r <= 16'b0101111011000111; rvalue_r <= 16'b0101111011011011;end
            11'b11001111111: begin lvalue_r <= 16'b0101111011011011; rvalue_r <= 16'b0101111011101110;end
            11'b11010000000: begin lvalue_r <= 16'b0101111011101110; rvalue_r <= 16'b0101111100000010;end
            11'b11010000001: begin lvalue_r <= 16'b0101111100000010; rvalue_r <= 16'b0101111100010101;end
            11'b11010000010: begin lvalue_r <= 16'b0101111100010101; rvalue_r <= 16'b0101111100101001;end
            11'b11010000011: begin lvalue_r <= 16'b0101111100101001; rvalue_r <= 16'b0101111100111100;end
            11'b11010000100: begin lvalue_r <= 16'b0101111100111100; rvalue_r <= 16'b0101111101010000;end
            11'b11010000101: begin lvalue_r <= 16'b0101111101010000; rvalue_r <= 16'b0101111101100011;end
            11'b11010000110: begin lvalue_r <= 16'b0101111101100011; rvalue_r <= 16'b0101111101110111;end
            11'b11010000111: begin lvalue_r <= 16'b0101111101110111; rvalue_r <= 16'b0101111110001011;end
            11'b11010001000: begin lvalue_r <= 16'b0101111110001011; rvalue_r <= 16'b0101111110011110;end
            11'b11010001001: begin lvalue_r <= 16'b0101111110011110; rvalue_r <= 16'b0101111110110010;end
            11'b11010001010: begin lvalue_r <= 16'b0101111110110010; rvalue_r <= 16'b0101111111000101;end
            11'b11010001011: begin lvalue_r <= 16'b0101111111000101; rvalue_r <= 16'b0101111111011001;end
            11'b11010001100: begin lvalue_r <= 16'b0101111111011001; rvalue_r <= 16'b0101111111101101;end
            11'b11010001101: begin lvalue_r <= 16'b0101111111101101; rvalue_r <= 16'b0110000000000000;end
            11'b11010001110: begin lvalue_r <= 16'b0110000000000000; rvalue_r <= 16'b0110000000010100;end
            11'b11010001111: begin lvalue_r <= 16'b0110000000010100; rvalue_r <= 16'b0110000000100111;end
            11'b11010010000: begin lvalue_r <= 16'b0110000000100111; rvalue_r <= 16'b0110000000111011;end
            11'b11010010001: begin lvalue_r <= 16'b0110000000111011; rvalue_r <= 16'b0110000001001111;end
            11'b11010010010: begin lvalue_r <= 16'b0110000001001111; rvalue_r <= 16'b0110000001100011;end
            11'b11010010011: begin lvalue_r <= 16'b0110000001100011; rvalue_r <= 16'b0110000001110110;end
            11'b11010010100: begin lvalue_r <= 16'b0110000001110110; rvalue_r <= 16'b0110000010001010;end
            11'b11010010101: begin lvalue_r <= 16'b0110000010001010; rvalue_r <= 16'b0110000010011110;end
            11'b11010010110: begin lvalue_r <= 16'b0110000010011110; rvalue_r <= 16'b0110000010110001;end
            11'b11010010111: begin lvalue_r <= 16'b0110000010110001; rvalue_r <= 16'b0110000011000101;end
            11'b11010011000: begin lvalue_r <= 16'b0110000011000101; rvalue_r <= 16'b0110000011011001;end
            11'b11010011001: begin lvalue_r <= 16'b0110000011011001; rvalue_r <= 16'b0110000011101101;end
            11'b11010011010: begin lvalue_r <= 16'b0110000011101101; rvalue_r <= 16'b0110000100000000;end
            11'b11010011011: begin lvalue_r <= 16'b0110000100000000; rvalue_r <= 16'b0110000100010100;end
            11'b11010011100: begin lvalue_r <= 16'b0110000100010100; rvalue_r <= 16'b0110000100101000;end
            11'b11010011101: begin lvalue_r <= 16'b0110000100101000; rvalue_r <= 16'b0110000100111100;end
            11'b11010011110: begin lvalue_r <= 16'b0110000100111100; rvalue_r <= 16'b0110000101010000;end
            11'b11010011111: begin lvalue_r <= 16'b0110000101010000; rvalue_r <= 16'b0110000101100011;end
            11'b11010100000: begin lvalue_r <= 16'b0110000101100011; rvalue_r <= 16'b0110000101110111;end
            11'b11010100001: begin lvalue_r <= 16'b0110000101110111; rvalue_r <= 16'b0110000110001011;end
            11'b11010100010: begin lvalue_r <= 16'b0110000110001011; rvalue_r <= 16'b0110000110011111;end
            11'b11010100011: begin lvalue_r <= 16'b0110000110011111; rvalue_r <= 16'b0110000110110011;end
            11'b11010100100: begin lvalue_r <= 16'b0110000110110011; rvalue_r <= 16'b0110000111000111;end
            11'b11010100101: begin lvalue_r <= 16'b0110000111000111; rvalue_r <= 16'b0110000111011011;end
            11'b11010100110: begin lvalue_r <= 16'b0110000111011011; rvalue_r <= 16'b0110000111101111;end
            11'b11010100111: begin lvalue_r <= 16'b0110000111101111; rvalue_r <= 16'b0110001000000011;end
            11'b11010101000: begin lvalue_r <= 16'b0110001000000011; rvalue_r <= 16'b0110001000010111;end
            11'b11010101001: begin lvalue_r <= 16'b0110001000010111; rvalue_r <= 16'b0110001000101010;end
            11'b11010101010: begin lvalue_r <= 16'b0110001000101010; rvalue_r <= 16'b0110001000111110;end
            11'b11010101011: begin lvalue_r <= 16'b0110001000111110; rvalue_r <= 16'b0110001001010010;end
            11'b11010101100: begin lvalue_r <= 16'b0110001001010010; rvalue_r <= 16'b0110001001100110;end
            11'b11010101101: begin lvalue_r <= 16'b0110001001100110; rvalue_r <= 16'b0110001001111010;end
            11'b11010101110: begin lvalue_r <= 16'b0110001001111010; rvalue_r <= 16'b0110001010001110;end
            11'b11010101111: begin lvalue_r <= 16'b0110001010001110; rvalue_r <= 16'b0110001010100010;end
            11'b11010110000: begin lvalue_r <= 16'b0110001010100010; rvalue_r <= 16'b0110001010110110;end
            11'b11010110001: begin lvalue_r <= 16'b0110001010110110; rvalue_r <= 16'b0110001011001011;end
            11'b11010110010: begin lvalue_r <= 16'b0110001011001011; rvalue_r <= 16'b0110001011011111;end
            11'b11010110011: begin lvalue_r <= 16'b0110001011011111; rvalue_r <= 16'b0110001011110011;end
            11'b11010110100: begin lvalue_r <= 16'b0110001011110011; rvalue_r <= 16'b0110001100000111;end
            11'b11010110101: begin lvalue_r <= 16'b0110001100000111; rvalue_r <= 16'b0110001100011011;end
            11'b11010110110: begin lvalue_r <= 16'b0110001100011011; rvalue_r <= 16'b0110001100101111;end
            11'b11010110111: begin lvalue_r <= 16'b0110001100101111; rvalue_r <= 16'b0110001101000011;end
            11'b11010111000: begin lvalue_r <= 16'b0110001101000011; rvalue_r <= 16'b0110001101010111;end
            11'b11010111001: begin lvalue_r <= 16'b0110001101010111; rvalue_r <= 16'b0110001101101011;end
            11'b11010111010: begin lvalue_r <= 16'b0110001101101011; rvalue_r <= 16'b0110001101111111;end
            11'b11010111011: begin lvalue_r <= 16'b0110001101111111; rvalue_r <= 16'b0110001110010100;end
            11'b11010111100: begin lvalue_r <= 16'b0110001110010100; rvalue_r <= 16'b0110001110101000;end
            11'b11010111101: begin lvalue_r <= 16'b0110001110101000; rvalue_r <= 16'b0110001110111100;end
            11'b11010111110: begin lvalue_r <= 16'b0110001110111100; rvalue_r <= 16'b0110001111010000;end
            11'b11010111111: begin lvalue_r <= 16'b0110001111010000; rvalue_r <= 16'b0110001111100100;end
            11'b11011000000: begin lvalue_r <= 16'b0110001111100100; rvalue_r <= 16'b0110001111111001;end
            11'b11011000001: begin lvalue_r <= 16'b0110001111111001; rvalue_r <= 16'b0110010000001101;end
            11'b11011000010: begin lvalue_r <= 16'b0110010000001101; rvalue_r <= 16'b0110010000100001;end
            11'b11011000011: begin lvalue_r <= 16'b0110010000100001; rvalue_r <= 16'b0110010000110101;end
            11'b11011000100: begin lvalue_r <= 16'b0110010000110101; rvalue_r <= 16'b0110010001001010;end
            11'b11011000101: begin lvalue_r <= 16'b0110010001001010; rvalue_r <= 16'b0110010001011110;end
            11'b11011000110: begin lvalue_r <= 16'b0110010001011110; rvalue_r <= 16'b0110010001110010;end
            11'b11011000111: begin lvalue_r <= 16'b0110010001110010; rvalue_r <= 16'b0110010010000111;end
            11'b11011001000: begin lvalue_r <= 16'b0110010010000111; rvalue_r <= 16'b0110010010011011;end
            11'b11011001001: begin lvalue_r <= 16'b0110010010011011; rvalue_r <= 16'b0110010010101111;end
            11'b11011001010: begin lvalue_r <= 16'b0110010010101111; rvalue_r <= 16'b0110010011000100;end
            11'b11011001011: begin lvalue_r <= 16'b0110010011000100; rvalue_r <= 16'b0110010011011000;end
            11'b11011001100: begin lvalue_r <= 16'b0110010011011000; rvalue_r <= 16'b0110010011101100;end
            11'b11011001101: begin lvalue_r <= 16'b0110010011101100; rvalue_r <= 16'b0110010100000001;end
            11'b11011001110: begin lvalue_r <= 16'b0110010100000001; rvalue_r <= 16'b0110010100010101;end
            11'b11011001111: begin lvalue_r <= 16'b0110010100010101; rvalue_r <= 16'b0110010100101001;end
            11'b11011010000: begin lvalue_r <= 16'b0110010100101001; rvalue_r <= 16'b0110010100111110;end
            11'b11011010001: begin lvalue_r <= 16'b0110010100111110; rvalue_r <= 16'b0110010101010010;end
            11'b11011010010: begin lvalue_r <= 16'b0110010101010010; rvalue_r <= 16'b0110010101100111;end
            11'b11011010011: begin lvalue_r <= 16'b0110010101100111; rvalue_r <= 16'b0110010101111011;end
            11'b11011010100: begin lvalue_r <= 16'b0110010101111011; rvalue_r <= 16'b0110010110010000;end
            11'b11011010101: begin lvalue_r <= 16'b0110010110010000; rvalue_r <= 16'b0110010110100100;end
            11'b11011010110: begin lvalue_r <= 16'b0110010110100100; rvalue_r <= 16'b0110010110111001;end
            11'b11011010111: begin lvalue_r <= 16'b0110010110111001; rvalue_r <= 16'b0110010111001101;end
            11'b11011011000: begin lvalue_r <= 16'b0110010111001101; rvalue_r <= 16'b0110010111100010;end
            11'b11011011001: begin lvalue_r <= 16'b0110010111100010; rvalue_r <= 16'b0110010111110110;end
            11'b11011011010: begin lvalue_r <= 16'b0110010111110110; rvalue_r <= 16'b0110011000001011;end
            11'b11011011011: begin lvalue_r <= 16'b0110011000001011; rvalue_r <= 16'b0110011000011111;end
            11'b11011011100: begin lvalue_r <= 16'b0110011000011111; rvalue_r <= 16'b0110011000110100;end
            11'b11011011101: begin lvalue_r <= 16'b0110011000110100; rvalue_r <= 16'b0110011001001001;end
            11'b11011011110: begin lvalue_r <= 16'b0110011001001001; rvalue_r <= 16'b0110011001011101;end
            11'b11011011111: begin lvalue_r <= 16'b0110011001011101; rvalue_r <= 16'b0110011001110010;end
            11'b11011100000: begin lvalue_r <= 16'b0110011001110010; rvalue_r <= 16'b0110011010000110;end
            11'b11011100001: begin lvalue_r <= 16'b0110011010000110; rvalue_r <= 16'b0110011010011011;end
            11'b11011100010: begin lvalue_r <= 16'b0110011010011011; rvalue_r <= 16'b0110011010110000;end
            11'b11011100011: begin lvalue_r <= 16'b0110011010110000; rvalue_r <= 16'b0110011011000100;end
            11'b11011100100: begin lvalue_r <= 16'b0110011011000100; rvalue_r <= 16'b0110011011011001;end
            11'b11011100101: begin lvalue_r <= 16'b0110011011011001; rvalue_r <= 16'b0110011011101110;end
            11'b11011100110: begin lvalue_r <= 16'b0110011011101110; rvalue_r <= 16'b0110011100000010;end
            11'b11011100111: begin lvalue_r <= 16'b0110011100000010; rvalue_r <= 16'b0110011100010111;end
            11'b11011101000: begin lvalue_r <= 16'b0110011100010111; rvalue_r <= 16'b0110011100101100;end
            11'b11011101001: begin lvalue_r <= 16'b0110011100101100; rvalue_r <= 16'b0110011101000001;end
            11'b11011101010: begin lvalue_r <= 16'b0110011101000001; rvalue_r <= 16'b0110011101010101;end
            11'b11011101011: begin lvalue_r <= 16'b0110011101010101; rvalue_r <= 16'b0110011101101010;end
            11'b11011101100: begin lvalue_r <= 16'b0110011101101010; rvalue_r <= 16'b0110011101111111;end
            11'b11011101101: begin lvalue_r <= 16'b0110011101111111; rvalue_r <= 16'b0110011110010100;end
            11'b11011101110: begin lvalue_r <= 16'b0110011110010100; rvalue_r <= 16'b0110011110101000;end
            11'b11011101111: begin lvalue_r <= 16'b0110011110101000; rvalue_r <= 16'b0110011110111101;end
            11'b11011110000: begin lvalue_r <= 16'b0110011110111101; rvalue_r <= 16'b0110011111010010;end
            11'b11011110001: begin lvalue_r <= 16'b0110011111010010; rvalue_r <= 16'b0110011111100111;end
            11'b11011110010: begin lvalue_r <= 16'b0110011111100111; rvalue_r <= 16'b0110011111111100;end
            11'b11011110011: begin lvalue_r <= 16'b0110011111111100; rvalue_r <= 16'b0110100000010001;end
            11'b11011110100: begin lvalue_r <= 16'b0110100000010001; rvalue_r <= 16'b0110100000100101;end
            11'b11011110101: begin lvalue_r <= 16'b0110100000100101; rvalue_r <= 16'b0110100000111010;end
            11'b11011110110: begin lvalue_r <= 16'b0110100000111010; rvalue_r <= 16'b0110100001001111;end
            11'b11011110111: begin lvalue_r <= 16'b0110100001001111; rvalue_r <= 16'b0110100001100100;end
            11'b11011111000: begin lvalue_r <= 16'b0110100001100100; rvalue_r <= 16'b0110100001111001;end
            11'b11011111001: begin lvalue_r <= 16'b0110100001111001; rvalue_r <= 16'b0110100010001110;end
            11'b11011111010: begin lvalue_r <= 16'b0110100010001110; rvalue_r <= 16'b0110100010100011;end
            11'b11011111011: begin lvalue_r <= 16'b0110100010100011; rvalue_r <= 16'b0110100010111000;end
            11'b11011111100: begin lvalue_r <= 16'b0110100010111000; rvalue_r <= 16'b0110100011001101;end
            11'b11011111101: begin lvalue_r <= 16'b0110100011001101; rvalue_r <= 16'b0110100011100010;end
            11'b11011111110: begin lvalue_r <= 16'b0110100011100010; rvalue_r <= 16'b0110100011110111;end
            11'b11011111111: begin lvalue_r <= 16'b0110100011110111; rvalue_r <= 16'b0110100100001100;end
            11'b11100000000: begin lvalue_r <= 16'b0110100100001100; rvalue_r <= 16'b0110100100100001;end
            11'b11100000001: begin lvalue_r <= 16'b0110100100100001; rvalue_r <= 16'b0110100100110110;end
            11'b11100000010: begin lvalue_r <= 16'b0110100100110110; rvalue_r <= 16'b0110100101001011;end
            11'b11100000011: begin lvalue_r <= 16'b0110100101001011; rvalue_r <= 16'b0110100101100000;end
            11'b11100000100: begin lvalue_r <= 16'b0110100101100000; rvalue_r <= 16'b0110100101110101;end
            11'b11100000101: begin lvalue_r <= 16'b0110100101110101; rvalue_r <= 16'b0110100110001010;end
            11'b11100000110: begin lvalue_r <= 16'b0110100110001010; rvalue_r <= 16'b0110100110100000;end
            11'b11100000111: begin lvalue_r <= 16'b0110100110100000; rvalue_r <= 16'b0110100110110101;end
            11'b11100001000: begin lvalue_r <= 16'b0110100110110101; rvalue_r <= 16'b0110100111001010;end
            11'b11100001001: begin lvalue_r <= 16'b0110100111001010; rvalue_r <= 16'b0110100111011111;end
            11'b11100001010: begin lvalue_r <= 16'b0110100111011111; rvalue_r <= 16'b0110100111110100;end
            11'b11100001011: begin lvalue_r <= 16'b0110100111110100; rvalue_r <= 16'b0110101000001001;end
            11'b11100001100: begin lvalue_r <= 16'b0110101000001001; rvalue_r <= 16'b0110101000011111;end
            11'b11100001101: begin lvalue_r <= 16'b0110101000011111; rvalue_r <= 16'b0110101000110100;end
            11'b11100001110: begin lvalue_r <= 16'b0110101000110100; rvalue_r <= 16'b0110101001001001;end
            11'b11100001111: begin lvalue_r <= 16'b0110101001001001; rvalue_r <= 16'b0110101001011110;end
            11'b11100010000: begin lvalue_r <= 16'b0110101001011110; rvalue_r <= 16'b0110101001110011;end
            11'b11100010001: begin lvalue_r <= 16'b0110101001110011; rvalue_r <= 16'b0110101010001001;end
            11'b11100010010: begin lvalue_r <= 16'b0110101010001001; rvalue_r <= 16'b0110101010011110;end
            11'b11100010011: begin lvalue_r <= 16'b0110101010011110; rvalue_r <= 16'b0110101010110011;end
            11'b11100010100: begin lvalue_r <= 16'b0110101010110011; rvalue_r <= 16'b0110101011001001;end
            11'b11100010101: begin lvalue_r <= 16'b0110101011001001; rvalue_r <= 16'b0110101011011110;end
            11'b11100010110: begin lvalue_r <= 16'b0110101011011110; rvalue_r <= 16'b0110101011110011;end
            11'b11100010111: begin lvalue_r <= 16'b0110101011110011; rvalue_r <= 16'b0110101100001001;end
            11'b11100011000: begin lvalue_r <= 16'b0110101100001001; rvalue_r <= 16'b0110101100011110;end
            11'b11100011001: begin lvalue_r <= 16'b0110101100011110; rvalue_r <= 16'b0110101100110011;end
            11'b11100011010: begin lvalue_r <= 16'b0110101100110011; rvalue_r <= 16'b0110101101001001;end
            11'b11100011011: begin lvalue_r <= 16'b0110101101001001; rvalue_r <= 16'b0110101101011110;end
            11'b11100011100: begin lvalue_r <= 16'b0110101101011110; rvalue_r <= 16'b0110101101110100;end
            11'b11100011101: begin lvalue_r <= 16'b0110101101110100; rvalue_r <= 16'b0110101110001001;end
            11'b11100011110: begin lvalue_r <= 16'b0110101110001001; rvalue_r <= 16'b0110101110011110;end
            11'b11100011111: begin lvalue_r <= 16'b0110101110011110; rvalue_r <= 16'b0110101110110100;end
            11'b11100100000: begin lvalue_r <= 16'b0110101110110100; rvalue_r <= 16'b0110101111001001;end
            11'b11100100001: begin lvalue_r <= 16'b0110101111001001; rvalue_r <= 16'b0110101111011111;end
            11'b11100100010: begin lvalue_r <= 16'b0110101111011111; rvalue_r <= 16'b0110101111110100;end
            11'b11100100011: begin lvalue_r <= 16'b0110101111110100; rvalue_r <= 16'b0110110000001010;end
            11'b11100100100: begin lvalue_r <= 16'b0110110000001010; rvalue_r <= 16'b0110110000011111;end
            11'b11100100101: begin lvalue_r <= 16'b0110110000011111; rvalue_r <= 16'b0110110000110101;end
            11'b11100100110: begin lvalue_r <= 16'b0110110000110101; rvalue_r <= 16'b0110110001001010;end
            11'b11100100111: begin lvalue_r <= 16'b0110110001001010; rvalue_r <= 16'b0110110001100000;end
            11'b11100101000: begin lvalue_r <= 16'b0110110001100000; rvalue_r <= 16'b0110110001110110;end
            11'b11100101001: begin lvalue_r <= 16'b0110110001110110; rvalue_r <= 16'b0110110010001011;end
            11'b11100101010: begin lvalue_r <= 16'b0110110010001011; rvalue_r <= 16'b0110110010100001;end
            11'b11100101011: begin lvalue_r <= 16'b0110110010100001; rvalue_r <= 16'b0110110010110110;end
            11'b11100101100: begin lvalue_r <= 16'b0110110010110110; rvalue_r <= 16'b0110110011001100;end
            11'b11100101101: begin lvalue_r <= 16'b0110110011001100; rvalue_r <= 16'b0110110011100010;end
            11'b11100101110: begin lvalue_r <= 16'b0110110011100010; rvalue_r <= 16'b0110110011110111;end
            11'b11100101111: begin lvalue_r <= 16'b0110110011110111; rvalue_r <= 16'b0110110100001101;end
            11'b11100110000: begin lvalue_r <= 16'b0110110100001101; rvalue_r <= 16'b0110110100100011;end
            11'b11100110001: begin lvalue_r <= 16'b0110110100100011; rvalue_r <= 16'b0110110100111000;end
            11'b11100110010: begin lvalue_r <= 16'b0110110100111000; rvalue_r <= 16'b0110110101001110;end
            11'b11100110011: begin lvalue_r <= 16'b0110110101001110; rvalue_r <= 16'b0110110101100100;end
            11'b11100110100: begin lvalue_r <= 16'b0110110101100100; rvalue_r <= 16'b0110110101111010;end
            11'b11100110101: begin lvalue_r <= 16'b0110110101111010; rvalue_r <= 16'b0110110110001111;end
            11'b11100110110: begin lvalue_r <= 16'b0110110110001111; rvalue_r <= 16'b0110110110100101;end
            11'b11100110111: begin lvalue_r <= 16'b0110110110100101; rvalue_r <= 16'b0110110110111011;end
            11'b11100111000: begin lvalue_r <= 16'b0110110110111011; rvalue_r <= 16'b0110110111010001;end
            11'b11100111001: begin lvalue_r <= 16'b0110110111010001; rvalue_r <= 16'b0110110111100111;end
            11'b11100111010: begin lvalue_r <= 16'b0110110111100111; rvalue_r <= 16'b0110110111111100;end
            11'b11100111011: begin lvalue_r <= 16'b0110110111111100; rvalue_r <= 16'b0110111000010010;end
            11'b11100111100: begin lvalue_r <= 16'b0110111000010010; rvalue_r <= 16'b0110111000101000;end
            11'b11100111101: begin lvalue_r <= 16'b0110111000101000; rvalue_r <= 16'b0110111000111110;end
            11'b11100111110: begin lvalue_r <= 16'b0110111000111110; rvalue_r <= 16'b0110111001010100;end
            11'b11100111111: begin lvalue_r <= 16'b0110111001010100; rvalue_r <= 16'b0110111001101010;end
            11'b11101000000: begin lvalue_r <= 16'b0110111001101010; rvalue_r <= 16'b0110111010000000;end
            11'b11101000001: begin lvalue_r <= 16'b0110111010000000; rvalue_r <= 16'b0110111010010110;end
            11'b11101000010: begin lvalue_r <= 16'b0110111010010110; rvalue_r <= 16'b0110111010101100;end
            11'b11101000011: begin lvalue_r <= 16'b0110111010101100; rvalue_r <= 16'b0110111011000010;end
            11'b11101000100: begin lvalue_r <= 16'b0110111011000010; rvalue_r <= 16'b0110111011011000;end
            11'b11101000101: begin lvalue_r <= 16'b0110111011011000; rvalue_r <= 16'b0110111011101110;end
            11'b11101000110: begin lvalue_r <= 16'b0110111011101110; rvalue_r <= 16'b0110111100000100;end
            11'b11101000111: begin lvalue_r <= 16'b0110111100000100; rvalue_r <= 16'b0110111100011010;end
            11'b11101001000: begin lvalue_r <= 16'b0110111100011010; rvalue_r <= 16'b0110111100110000;end
            11'b11101001001: begin lvalue_r <= 16'b0110111100110000; rvalue_r <= 16'b0110111101000110;end
            11'b11101001010: begin lvalue_r <= 16'b0110111101000110; rvalue_r <= 16'b0110111101011100;end
            11'b11101001011: begin lvalue_r <= 16'b0110111101011100; rvalue_r <= 16'b0110111101110010;end
            11'b11101001100: begin lvalue_r <= 16'b0110111101110010; rvalue_r <= 16'b0110111110001000;end
            11'b11101001101: begin lvalue_r <= 16'b0110111110001000; rvalue_r <= 16'b0110111110011110;end
            11'b11101001110: begin lvalue_r <= 16'b0110111110011110; rvalue_r <= 16'b0110111110110100;end
            11'b11101001111: begin lvalue_r <= 16'b0110111110110100; rvalue_r <= 16'b0110111111001010;end
            11'b11101010000: begin lvalue_r <= 16'b0110111111001010; rvalue_r <= 16'b0110111111100001;end
            11'b11101010001: begin lvalue_r <= 16'b0110111111100001; rvalue_r <= 16'b0110111111110111;end
            11'b11101010010: begin lvalue_r <= 16'b0110111111110111; rvalue_r <= 16'b0111000000001101;end
            11'b11101010011: begin lvalue_r <= 16'b0111000000001101; rvalue_r <= 16'b0111000000100011;end
            11'b11101010100: begin lvalue_r <= 16'b0111000000100011; rvalue_r <= 16'b0111000000111001;end
            11'b11101010101: begin lvalue_r <= 16'b0111000000111001; rvalue_r <= 16'b0111000001010000;end
            11'b11101010110: begin lvalue_r <= 16'b0111000001010000; rvalue_r <= 16'b0111000001100110;end
            11'b11101010111: begin lvalue_r <= 16'b0111000001100110; rvalue_r <= 16'b0111000001111100;end
            11'b11101011000: begin lvalue_r <= 16'b0111000001111100; rvalue_r <= 16'b0111000010010010;end
            11'b11101011001: begin lvalue_r <= 16'b0111000010010010; rvalue_r <= 16'b0111000010101001;end
            11'b11101011010: begin lvalue_r <= 16'b0111000010101001; rvalue_r <= 16'b0111000010111111;end
            11'b11101011011: begin lvalue_r <= 16'b0111000010111111; rvalue_r <= 16'b0111000011010101;end
            11'b11101011100: begin lvalue_r <= 16'b0111000011010101; rvalue_r <= 16'b0111000011101100;end
            11'b11101011101: begin lvalue_r <= 16'b0111000011101100; rvalue_r <= 16'b0111000100000010;end
            11'b11101011110: begin lvalue_r <= 16'b0111000100000010; rvalue_r <= 16'b0111000100011000;end
            11'b11101011111: begin lvalue_r <= 16'b0111000100011000; rvalue_r <= 16'b0111000100101111;end
            11'b11101100000: begin lvalue_r <= 16'b0111000100101111; rvalue_r <= 16'b0111000101000101;end
            11'b11101100001: begin lvalue_r <= 16'b0111000101000101; rvalue_r <= 16'b0111000101011100;end
            11'b11101100010: begin lvalue_r <= 16'b0111000101011100; rvalue_r <= 16'b0111000101110010;end
            11'b11101100011: begin lvalue_r <= 16'b0111000101110010; rvalue_r <= 16'b0111000110001000;end
            11'b11101100100: begin lvalue_r <= 16'b0111000110001000; rvalue_r <= 16'b0111000110011111;end
            11'b11101100101: begin lvalue_r <= 16'b0111000110011111; rvalue_r <= 16'b0111000110110101;end
            11'b11101100110: begin lvalue_r <= 16'b0111000110110101; rvalue_r <= 16'b0111000111001100;end
            11'b11101100111: begin lvalue_r <= 16'b0111000111001100; rvalue_r <= 16'b0111000111100010;end
            11'b11101101000: begin lvalue_r <= 16'b0111000111100010; rvalue_r <= 16'b0111000111111001;end
            11'b11101101001: begin lvalue_r <= 16'b0111000111111001; rvalue_r <= 16'b0111001000001111;end
            11'b11101101010: begin lvalue_r <= 16'b0111001000001111; rvalue_r <= 16'b0111001000100110;end
            11'b11101101011: begin lvalue_r <= 16'b0111001000100110; rvalue_r <= 16'b0111001000111101;end
            11'b11101101100: begin lvalue_r <= 16'b0111001000111101; rvalue_r <= 16'b0111001001010011;end
            11'b11101101101: begin lvalue_r <= 16'b0111001001010011; rvalue_r <= 16'b0111001001101010;end
            11'b11101101110: begin lvalue_r <= 16'b0111001001101010; rvalue_r <= 16'b0111001010000000;end
            11'b11101101111: begin lvalue_r <= 16'b0111001010000000; rvalue_r <= 16'b0111001010010111;end
            11'b11101110000: begin lvalue_r <= 16'b0111001010010111; rvalue_r <= 16'b0111001010101110;end
            11'b11101110001: begin lvalue_r <= 16'b0111001010101110; rvalue_r <= 16'b0111001011000100;end
            11'b11101110010: begin lvalue_r <= 16'b0111001011000100; rvalue_r <= 16'b0111001011011011;end
            11'b11101110011: begin lvalue_r <= 16'b0111001011011011; rvalue_r <= 16'b0111001011110010;end
            11'b11101110100: begin lvalue_r <= 16'b0111001011110010; rvalue_r <= 16'b0111001100001000;end
            11'b11101110101: begin lvalue_r <= 16'b0111001100001000; rvalue_r <= 16'b0111001100011111;end
            11'b11101110110: begin lvalue_r <= 16'b0111001100011111; rvalue_r <= 16'b0111001100110110;end
            11'b11101110111: begin lvalue_r <= 16'b0111001100110110; rvalue_r <= 16'b0111001101001101;end
            11'b11101111000: begin lvalue_r <= 16'b0111001101001101; rvalue_r <= 16'b0111001101100011;end
            11'b11101111001: begin lvalue_r <= 16'b0111001101100011; rvalue_r <= 16'b0111001101111010;end
            11'b11101111010: begin lvalue_r <= 16'b0111001101111010; rvalue_r <= 16'b0111001110010001;end
            11'b11101111011: begin lvalue_r <= 16'b0111001110010001; rvalue_r <= 16'b0111001110101000;end
            11'b11101111100: begin lvalue_r <= 16'b0111001110101000; rvalue_r <= 16'b0111001110111111;end
            11'b11101111101: begin lvalue_r <= 16'b0111001110111111; rvalue_r <= 16'b0111001111010101;end
            11'b11101111110: begin lvalue_r <= 16'b0111001111010101; rvalue_r <= 16'b0111001111101100;end
            11'b11101111111: begin lvalue_r <= 16'b0111001111101100; rvalue_r <= 16'b0111010000000011;end
            11'b11110000000: begin lvalue_r <= 16'b0111010000000011; rvalue_r <= 16'b0111010000011010;end
            11'b11110000001: begin lvalue_r <= 16'b0111010000011010; rvalue_r <= 16'b0111010000110001;end
            11'b11110000010: begin lvalue_r <= 16'b0111010000110001; rvalue_r <= 16'b0111010001001000;end
            11'b11110000011: begin lvalue_r <= 16'b0111010001001000; rvalue_r <= 16'b0111010001011111;end
            11'b11110000100: begin lvalue_r <= 16'b0111010001011111; rvalue_r <= 16'b0111010001110110;end
            11'b11110000101: begin lvalue_r <= 16'b0111010001110110; rvalue_r <= 16'b0111010010001101;end
            11'b11110000110: begin lvalue_r <= 16'b0111010010001101; rvalue_r <= 16'b0111010010100100;end
            11'b11110000111: begin lvalue_r <= 16'b0111010010100100; rvalue_r <= 16'b0111010010111011;end
            11'b11110001000: begin lvalue_r <= 16'b0111010010111011; rvalue_r <= 16'b0111010011010010;end
            11'b11110001001: begin lvalue_r <= 16'b0111010011010010; rvalue_r <= 16'b0111010011101001;end
            11'b11110001010: begin lvalue_r <= 16'b0111010011101001; rvalue_r <= 16'b0111010100000000;end
            11'b11110001011: begin lvalue_r <= 16'b0111010100000000; rvalue_r <= 16'b0111010100010111;end
            11'b11110001100: begin lvalue_r <= 16'b0111010100010111; rvalue_r <= 16'b0111010100101110;end
            11'b11110001101: begin lvalue_r <= 16'b0111010100101110; rvalue_r <= 16'b0111010101000101;end
            11'b11110001110: begin lvalue_r <= 16'b0111010101000101; rvalue_r <= 16'b0111010101011100;end
            11'b11110001111: begin lvalue_r <= 16'b0111010101011100; rvalue_r <= 16'b0111010101110011;end
            11'b11110010000: begin lvalue_r <= 16'b0111010101110011; rvalue_r <= 16'b0111010110001011;end
            11'b11110010001: begin lvalue_r <= 16'b0111010110001011; rvalue_r <= 16'b0111010110100010;end
            11'b11110010010: begin lvalue_r <= 16'b0111010110100010; rvalue_r <= 16'b0111010110111001;end
            11'b11110010011: begin lvalue_r <= 16'b0111010110111001; rvalue_r <= 16'b0111010111010000;end
            11'b11110010100: begin lvalue_r <= 16'b0111010111010000; rvalue_r <= 16'b0111010111100111;end
            11'b11110010101: begin lvalue_r <= 16'b0111010111100111; rvalue_r <= 16'b0111010111111111;end
            11'b11110010110: begin lvalue_r <= 16'b0111010111111111; rvalue_r <= 16'b0111011000010110;end
            11'b11110010111: begin lvalue_r <= 16'b0111011000010110; rvalue_r <= 16'b0111011000101101;end
            11'b11110011000: begin lvalue_r <= 16'b0111011000101101; rvalue_r <= 16'b0111011001000100;end
            11'b11110011001: begin lvalue_r <= 16'b0111011001000100; rvalue_r <= 16'b0111011001011100;end
            11'b11110011010: begin lvalue_r <= 16'b0111011001011100; rvalue_r <= 16'b0111011001110011;end
            11'b11110011011: begin lvalue_r <= 16'b0111011001110011; rvalue_r <= 16'b0111011010001010;end
            11'b11110011100: begin lvalue_r <= 16'b0111011010001010; rvalue_r <= 16'b0111011010100010;end
            11'b11110011101: begin lvalue_r <= 16'b0111011010100010; rvalue_r <= 16'b0111011010111001;end
            11'b11110011110: begin lvalue_r <= 16'b0111011010111001; rvalue_r <= 16'b0111011011010001;end
            11'b11110011111: begin lvalue_r <= 16'b0111011011010001; rvalue_r <= 16'b0111011011101000;end
            11'b11110100000: begin lvalue_r <= 16'b0111011011101000; rvalue_r <= 16'b0111011011111111;end
            11'b11110100001: begin lvalue_r <= 16'b0111011011111111; rvalue_r <= 16'b0111011100010111;end
            11'b11110100010: begin lvalue_r <= 16'b0111011100010111; rvalue_r <= 16'b0111011100101110;end
            11'b11110100011: begin lvalue_r <= 16'b0111011100101110; rvalue_r <= 16'b0111011101000110;end
            11'b11110100100: begin lvalue_r <= 16'b0111011101000110; rvalue_r <= 16'b0111011101011101;end
            11'b11110100101: begin lvalue_r <= 16'b0111011101011101; rvalue_r <= 16'b0111011101110101;end
            11'b11110100110: begin lvalue_r <= 16'b0111011101110101; rvalue_r <= 16'b0111011110001100;end
            11'b11110100111: begin lvalue_r <= 16'b0111011110001100; rvalue_r <= 16'b0111011110100100;end
            11'b11110101000: begin lvalue_r <= 16'b0111011110100100; rvalue_r <= 16'b0111011110111011;end
            11'b11110101001: begin lvalue_r <= 16'b0111011110111011; rvalue_r <= 16'b0111011111010011;end
            11'b11110101010: begin lvalue_r <= 16'b0111011111010011; rvalue_r <= 16'b0111011111101010;end
            11'b11110101011: begin lvalue_r <= 16'b0111011111101010; rvalue_r <= 16'b0111100000000010;end
            11'b11110101100: begin lvalue_r <= 16'b0111100000000010; rvalue_r <= 16'b0111100000011010;end
            11'b11110101101: begin lvalue_r <= 16'b0111100000011010; rvalue_r <= 16'b0111100000110001;end
            11'b11110101110: begin lvalue_r <= 16'b0111100000110001; rvalue_r <= 16'b0111100001001001;end
            11'b11110101111: begin lvalue_r <= 16'b0111100001001001; rvalue_r <= 16'b0111100001100001;end
            11'b11110110000: begin lvalue_r <= 16'b0111100001100001; rvalue_r <= 16'b0111100001111000;end
            11'b11110110001: begin lvalue_r <= 16'b0111100001111000; rvalue_r <= 16'b0111100010010000;end
            11'b11110110010: begin lvalue_r <= 16'b0111100010010000; rvalue_r <= 16'b0111100010101000;end
            11'b11110110011: begin lvalue_r <= 16'b0111100010101000; rvalue_r <= 16'b0111100010111111;end
            11'b11110110100: begin lvalue_r <= 16'b0111100010111111; rvalue_r <= 16'b0111100011010111;end
            11'b11110110101: begin lvalue_r <= 16'b0111100011010111; rvalue_r <= 16'b0111100011101111;end
            11'b11110110110: begin lvalue_r <= 16'b0111100011101111; rvalue_r <= 16'b0111100100000111;end
            11'b11110110111: begin lvalue_r <= 16'b0111100100000111; rvalue_r <= 16'b0111100100011111;end
            11'b11110111000: begin lvalue_r <= 16'b0111100100011111; rvalue_r <= 16'b0111100100110110;end
            11'b11110111001: begin lvalue_r <= 16'b0111100100110110; rvalue_r <= 16'b0111100101001110;end
            11'b11110111010: begin lvalue_r <= 16'b0111100101001110; rvalue_r <= 16'b0111100101100110;end
            11'b11110111011: begin lvalue_r <= 16'b0111100101100110; rvalue_r <= 16'b0111100101111110;end
            11'b11110111100: begin lvalue_r <= 16'b0111100101111110; rvalue_r <= 16'b0111100110010110;end
            11'b11110111101: begin lvalue_r <= 16'b0111100110010110; rvalue_r <= 16'b0111100110101110;end
            11'b11110111110: begin lvalue_r <= 16'b0111100110101110; rvalue_r <= 16'b0111100111000110;end
            11'b11110111111: begin lvalue_r <= 16'b0111100111000110; rvalue_r <= 16'b0111100111011110;end
            11'b11111000000: begin lvalue_r <= 16'b0111100111011110; rvalue_r <= 16'b0111100111110110;end
            11'b11111000001: begin lvalue_r <= 16'b0111100111110110; rvalue_r <= 16'b0111101000001110;end
            11'b11111000010: begin lvalue_r <= 16'b0111101000001110; rvalue_r <= 16'b0111101000100110;end
            11'b11111000011: begin lvalue_r <= 16'b0111101000100110; rvalue_r <= 16'b0111101000111110;end
            11'b11111000100: begin lvalue_r <= 16'b0111101000111110; rvalue_r <= 16'b0111101001010110;end
            11'b11111000101: begin lvalue_r <= 16'b0111101001010110; rvalue_r <= 16'b0111101001101110;end
            11'b11111000110: begin lvalue_r <= 16'b0111101001101110; rvalue_r <= 16'b0111101010000110;end
            11'b11111000111: begin lvalue_r <= 16'b0111101010000110; rvalue_r <= 16'b0111101010011110;end
            11'b11111001000: begin lvalue_r <= 16'b0111101010011110; rvalue_r <= 16'b0111101010110110;end
            11'b11111001001: begin lvalue_r <= 16'b0111101010110110; rvalue_r <= 16'b0111101011001110;end
            11'b11111001010: begin lvalue_r <= 16'b0111101011001110; rvalue_r <= 16'b0111101011100110;end
            11'b11111001011: begin lvalue_r <= 16'b0111101011100110; rvalue_r <= 16'b0111101011111110;end
            11'b11111001100: begin lvalue_r <= 16'b0111101011111110; rvalue_r <= 16'b0111101100010111;end
            11'b11111001101: begin lvalue_r <= 16'b0111101100010111; rvalue_r <= 16'b0111101100101111;end
            11'b11111001110: begin lvalue_r <= 16'b0111101100101111; rvalue_r <= 16'b0111101101000111;end
            11'b11111001111: begin lvalue_r <= 16'b0111101101000111; rvalue_r <= 16'b0111101101011111;end
            11'b11111010000: begin lvalue_r <= 16'b0111101101011111; rvalue_r <= 16'b0111101101111000;end
            11'b11111010001: begin lvalue_r <= 16'b0111101101111000; rvalue_r <= 16'b0111101110010000;end
            11'b11111010010: begin lvalue_r <= 16'b0111101110010000; rvalue_r <= 16'b0111101110101000;end
            11'b11111010011: begin lvalue_r <= 16'b0111101110101000; rvalue_r <= 16'b0111101111000000;end
            11'b11111010100: begin lvalue_r <= 16'b0111101111000000; rvalue_r <= 16'b0111101111011001;end
            11'b11111010101: begin lvalue_r <= 16'b0111101111011001; rvalue_r <= 16'b0111101111110001;end
            11'b11111010110: begin lvalue_r <= 16'b0111101111110001; rvalue_r <= 16'b0111110000001001;end
            11'b11111010111: begin lvalue_r <= 16'b0111110000001001; rvalue_r <= 16'b0111110000100010;end
            11'b11111011000: begin lvalue_r <= 16'b0111110000100010; rvalue_r <= 16'b0111110000111010;end
            11'b11111011001: begin lvalue_r <= 16'b0111110000111010; rvalue_r <= 16'b0111110001010011;end
            11'b11111011010: begin lvalue_r <= 16'b0111110001010011; rvalue_r <= 16'b0111110001101011;end
            11'b11111011011: begin lvalue_r <= 16'b0111110001101011; rvalue_r <= 16'b0111110010000011;end
            11'b11111011100: begin lvalue_r <= 16'b0111110010000011; rvalue_r <= 16'b0111110010011100;end
            11'b11111011101: begin lvalue_r <= 16'b0111110010011100; rvalue_r <= 16'b0111110010110100;end
            11'b11111011110: begin lvalue_r <= 16'b0111110010110100; rvalue_r <= 16'b0111110011001101;end
            11'b11111011111: begin lvalue_r <= 16'b0111110011001101; rvalue_r <= 16'b0111110011100101;end
            11'b11111100000: begin lvalue_r <= 16'b0111110011100101; rvalue_r <= 16'b0111110011111110;end
            11'b11111100001: begin lvalue_r <= 16'b0111110011111110; rvalue_r <= 16'b0111110100010111;end
            11'b11111100010: begin lvalue_r <= 16'b0111110100010111; rvalue_r <= 16'b0111110100101111;end
            11'b11111100011: begin lvalue_r <= 16'b0111110100101111; rvalue_r <= 16'b0111110101001000;end
            11'b11111100100: begin lvalue_r <= 16'b0111110101001000; rvalue_r <= 16'b0111110101100000;end
            11'b11111100101: begin lvalue_r <= 16'b0111110101100000; rvalue_r <= 16'b0111110101111001;end
            11'b11111100110: begin lvalue_r <= 16'b0111110101111001; rvalue_r <= 16'b0111110110010010;end
            11'b11111100111: begin lvalue_r <= 16'b0111110110010010; rvalue_r <= 16'b0111110110101010;end
            11'b11111101000: begin lvalue_r <= 16'b0111110110101010; rvalue_r <= 16'b0111110111000011;end
            11'b11111101001: begin lvalue_r <= 16'b0111110111000011; rvalue_r <= 16'b0111110111011100;end
            11'b11111101010: begin lvalue_r <= 16'b0111110111011100; rvalue_r <= 16'b0111110111110100;end
            11'b11111101011: begin lvalue_r <= 16'b0111110111110100; rvalue_r <= 16'b0111111000001101;end
            11'b11111101100: begin lvalue_r <= 16'b0111111000001101; rvalue_r <= 16'b0111111000100110;end
            11'b11111101101: begin lvalue_r <= 16'b0111111000100110; rvalue_r <= 16'b0111111000111111;end
            11'b11111101110: begin lvalue_r <= 16'b0111111000111111; rvalue_r <= 16'b0111111001011000;end
            11'b11111101111: begin lvalue_r <= 16'b0111111001011000; rvalue_r <= 16'b0111111001110000;end
            11'b11111110000: begin lvalue_r <= 16'b0111111001110000; rvalue_r <= 16'b0111111010001001;end
            11'b11111110001: begin lvalue_r <= 16'b0111111010001001; rvalue_r <= 16'b0111111010100010;end
            11'b11111110010: begin lvalue_r <= 16'b0111111010100010; rvalue_r <= 16'b0111111010111011;end
            11'b11111110011: begin lvalue_r <= 16'b0111111010111011; rvalue_r <= 16'b0111111011010100;end
            11'b11111110100: begin lvalue_r <= 16'b0111111011010100; rvalue_r <= 16'b0111111011101101;end
            11'b11111110101: begin lvalue_r <= 16'b0111111011101101; rvalue_r <= 16'b0111111100000110;end
            11'b11111110110: begin lvalue_r <= 16'b0111111100000110; rvalue_r <= 16'b0111111100011111;end
            11'b11111110111: begin lvalue_r <= 16'b0111111100011111; rvalue_r <= 16'b0111111100111000;end
            11'b11111111000: begin lvalue_r <= 16'b0111111100111000; rvalue_r <= 16'b0111111101010001;end
            11'b11111111001: begin lvalue_r <= 16'b0111111101010001; rvalue_r <= 16'b0111111101101010;end
            11'b11111111010: begin lvalue_r <= 16'b0111111101101010; rvalue_r <= 16'b0111111110000011;end
            11'b11111111011: begin lvalue_r <= 16'b0111111110000011; rvalue_r <= 16'b0111111110011100;end
            11'b11111111100: begin lvalue_r <= 16'b0111111110011100; rvalue_r <= 16'b0111111110110101;end
            11'b11111111101: begin lvalue_r <= 16'b0111111110110101; rvalue_r <= 16'b0111111111001110;end
            11'b11111111110: begin lvalue_r <= 16'b0111111111001110; rvalue_r <= 16'b0111111111100111;end
            11'b11111111111: begin lvalue_r <= 16'b0111111111100111; rvalue_r <= 16'b1000000000000000;end
            default: begin lvalue_r <= 16'b1111111111111111; rvalue_r <= 16'b1111111111111111;end
        endcase
        if(theta[0] == 1'b0)
            even <= 1'b1;
        else
            even <= 1'b0;
    end
    always @(posedge clk) begin
        if(even == 1'b1)
            out <= #1 lvalue_r;
        else
            out <= #1 ({1'b0,lvalue_r} + {1'b0,rvalue_r}) >> 1;
    end
endmodule